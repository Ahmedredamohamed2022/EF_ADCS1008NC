magic
tech sky130A
magscale 1 2
timestamp 1699926577
<< pwell >>
rect -1018 -298 1018 298
<< mvnmos >>
rect -800 -50 800 50
<< mvndiff >>
rect -858 17 -800 50
rect -858 -17 -846 17
rect -812 -17 -800 17
rect -858 -50 -800 -17
rect 800 17 858 50
rect 800 -17 812 17
rect 846 -17 858 17
rect 800 -50 858 -17
<< mvndiffc >>
rect -846 -17 -812 17
rect 812 -17 846 17
<< mvpsubdiff >>
rect -992 260 992 272
rect -992 226 -867 260
rect -833 226 -799 260
rect -765 226 -731 260
rect -697 226 -663 260
rect -629 226 -595 260
rect -561 226 -527 260
rect -493 226 -459 260
rect -425 226 -391 260
rect -357 226 -323 260
rect -289 226 -255 260
rect -221 226 -187 260
rect -153 226 -119 260
rect -85 226 -51 260
rect -17 226 17 260
rect 51 226 85 260
rect 119 226 153 260
rect 187 226 221 260
rect 255 226 289 260
rect 323 226 357 260
rect 391 226 425 260
rect 459 226 493 260
rect 527 226 561 260
rect 595 226 629 260
rect 663 226 697 260
rect 731 226 765 260
rect 799 226 833 260
rect 867 226 992 260
rect -992 214 992 226
rect -992 153 -934 214
rect -992 119 -980 153
rect -946 119 -934 153
rect 934 153 992 214
rect -992 85 -934 119
rect -992 51 -980 85
rect -946 51 -934 85
rect -992 17 -934 51
rect 934 119 946 153
rect 980 119 992 153
rect 934 85 992 119
rect 934 51 946 85
rect 980 51 992 85
rect -992 -17 -980 17
rect -946 -17 -934 17
rect -992 -51 -934 -17
rect 934 17 992 51
rect 934 -17 946 17
rect 980 -17 992 17
rect -992 -85 -980 -51
rect -946 -85 -934 -51
rect -992 -119 -934 -85
rect -992 -153 -980 -119
rect -946 -153 -934 -119
rect 934 -51 992 -17
rect 934 -85 946 -51
rect 980 -85 992 -51
rect 934 -119 992 -85
rect -992 -214 -934 -153
rect 934 -153 946 -119
rect 980 -153 992 -119
rect 934 -214 992 -153
rect -992 -226 992 -214
rect -992 -260 -867 -226
rect -833 -260 -799 -226
rect -765 -260 -731 -226
rect -697 -260 -663 -226
rect -629 -260 -595 -226
rect -561 -260 -527 -226
rect -493 -260 -459 -226
rect -425 -260 -391 -226
rect -357 -260 -323 -226
rect -289 -260 -255 -226
rect -221 -260 -187 -226
rect -153 -260 -119 -226
rect -85 -260 -51 -226
rect -17 -260 17 -226
rect 51 -260 85 -226
rect 119 -260 153 -226
rect 187 -260 221 -226
rect 255 -260 289 -226
rect 323 -260 357 -226
rect 391 -260 425 -226
rect 459 -260 493 -226
rect 527 -260 561 -226
rect 595 -260 629 -226
rect 663 -260 697 -226
rect 731 -260 765 -226
rect 799 -260 833 -226
rect 867 -260 992 -226
rect -992 -272 992 -260
<< mvpsubdiffcont >>
rect -867 226 -833 260
rect -799 226 -765 260
rect -731 226 -697 260
rect -663 226 -629 260
rect -595 226 -561 260
rect -527 226 -493 260
rect -459 226 -425 260
rect -391 226 -357 260
rect -323 226 -289 260
rect -255 226 -221 260
rect -187 226 -153 260
rect -119 226 -85 260
rect -51 226 -17 260
rect 17 226 51 260
rect 85 226 119 260
rect 153 226 187 260
rect 221 226 255 260
rect 289 226 323 260
rect 357 226 391 260
rect 425 226 459 260
rect 493 226 527 260
rect 561 226 595 260
rect 629 226 663 260
rect 697 226 731 260
rect 765 226 799 260
rect 833 226 867 260
rect -980 119 -946 153
rect -980 51 -946 85
rect 946 119 980 153
rect 946 51 980 85
rect -980 -17 -946 17
rect 946 -17 980 17
rect -980 -85 -946 -51
rect -980 -153 -946 -119
rect 946 -85 980 -51
rect 946 -153 980 -119
rect -867 -260 -833 -226
rect -799 -260 -765 -226
rect -731 -260 -697 -226
rect -663 -260 -629 -226
rect -595 -260 -561 -226
rect -527 -260 -493 -226
rect -459 -260 -425 -226
rect -391 -260 -357 -226
rect -323 -260 -289 -226
rect -255 -260 -221 -226
rect -187 -260 -153 -226
rect -119 -260 -85 -226
rect -51 -260 -17 -226
rect 17 -260 51 -226
rect 85 -260 119 -226
rect 153 -260 187 -226
rect 221 -260 255 -226
rect 289 -260 323 -226
rect 357 -260 391 -226
rect 425 -260 459 -226
rect 493 -260 527 -226
rect 561 -260 595 -226
rect 629 -260 663 -226
rect 697 -260 731 -226
rect 765 -260 799 -226
rect 833 -260 867 -226
<< poly >>
rect -800 122 800 138
rect -800 88 -765 122
rect -731 88 -697 122
rect -663 88 -629 122
rect -595 88 -561 122
rect -527 88 -493 122
rect -459 88 -425 122
rect -391 88 -357 122
rect -323 88 -289 122
rect -255 88 -221 122
rect -187 88 -153 122
rect -119 88 -85 122
rect -51 88 -17 122
rect 17 88 51 122
rect 85 88 119 122
rect 153 88 187 122
rect 221 88 255 122
rect 289 88 323 122
rect 357 88 391 122
rect 425 88 459 122
rect 493 88 527 122
rect 561 88 595 122
rect 629 88 663 122
rect 697 88 731 122
rect 765 88 800 122
rect -800 50 800 88
rect -800 -88 800 -50
rect -800 -122 -765 -88
rect -731 -122 -697 -88
rect -663 -122 -629 -88
rect -595 -122 -561 -88
rect -527 -122 -493 -88
rect -459 -122 -425 -88
rect -391 -122 -357 -88
rect -323 -122 -289 -88
rect -255 -122 -221 -88
rect -187 -122 -153 -88
rect -119 -122 -85 -88
rect -51 -122 -17 -88
rect 17 -122 51 -88
rect 85 -122 119 -88
rect 153 -122 187 -88
rect 221 -122 255 -88
rect 289 -122 323 -88
rect 357 -122 391 -88
rect 425 -122 459 -88
rect 493 -122 527 -88
rect 561 -122 595 -88
rect 629 -122 663 -88
rect 697 -122 731 -88
rect 765 -122 800 -88
rect -800 -138 800 -122
<< polycont >>
rect -765 88 -731 122
rect -697 88 -663 122
rect -629 88 -595 122
rect -561 88 -527 122
rect -493 88 -459 122
rect -425 88 -391 122
rect -357 88 -323 122
rect -289 88 -255 122
rect -221 88 -187 122
rect -153 88 -119 122
rect -85 88 -51 122
rect -17 88 17 122
rect 51 88 85 122
rect 119 88 153 122
rect 187 88 221 122
rect 255 88 289 122
rect 323 88 357 122
rect 391 88 425 122
rect 459 88 493 122
rect 527 88 561 122
rect 595 88 629 122
rect 663 88 697 122
rect 731 88 765 122
rect -765 -122 -731 -88
rect -697 -122 -663 -88
rect -629 -122 -595 -88
rect -561 -122 -527 -88
rect -493 -122 -459 -88
rect -425 -122 -391 -88
rect -357 -122 -323 -88
rect -289 -122 -255 -88
rect -221 -122 -187 -88
rect -153 -122 -119 -88
rect -85 -122 -51 -88
rect -17 -122 17 -88
rect 51 -122 85 -88
rect 119 -122 153 -88
rect 187 -122 221 -88
rect 255 -122 289 -88
rect 323 -122 357 -88
rect 391 -122 425 -88
rect 459 -122 493 -88
rect 527 -122 561 -88
rect 595 -122 629 -88
rect 663 -122 697 -88
rect 731 -122 765 -88
<< locali >>
rect -980 226 -917 260
rect -883 226 -867 260
rect -811 226 -799 260
rect -739 226 -731 260
rect -667 226 -663 260
rect -561 226 -557 260
rect -493 226 -485 260
rect -425 226 -413 260
rect -357 226 -341 260
rect -289 226 -269 260
rect -221 226 -197 260
rect -153 226 -125 260
rect -85 226 -53 260
rect -17 226 17 260
rect 53 226 85 260
rect 125 226 153 260
rect 197 226 221 260
rect 269 226 289 260
rect 341 226 357 260
rect 413 226 425 260
rect 485 226 493 260
rect 557 226 561 260
rect 663 226 667 260
rect 731 226 739 260
rect 799 226 811 260
rect 867 226 883 260
rect 917 226 980 260
rect -980 153 -946 226
rect 946 153 980 226
rect -980 85 -946 119
rect -800 88 -773 122
rect -731 88 -701 122
rect -663 88 -629 122
rect -595 88 -561 122
rect -523 88 -493 122
rect -451 88 -425 122
rect -379 88 -357 122
rect -307 88 -289 122
rect -235 88 -221 122
rect -163 88 -153 122
rect -91 88 -85 122
rect -19 88 -17 122
rect 17 88 19 122
rect 85 88 91 122
rect 153 88 163 122
rect 221 88 235 122
rect 289 88 307 122
rect 357 88 379 122
rect 425 88 451 122
rect 493 88 523 122
rect 561 88 595 122
rect 629 88 663 122
rect 701 88 731 122
rect 773 88 800 122
rect 946 85 980 119
rect -980 17 -946 51
rect -980 -51 -946 -17
rect -846 17 -812 54
rect -846 -54 -812 -17
rect 812 17 846 54
rect 812 -54 846 -17
rect 946 17 980 51
rect 946 -51 980 -17
rect -980 -119 -946 -85
rect -800 -122 -773 -88
rect -731 -122 -701 -88
rect -663 -122 -629 -88
rect -595 -122 -561 -88
rect -523 -122 -493 -88
rect -451 -122 -425 -88
rect -379 -122 -357 -88
rect -307 -122 -289 -88
rect -235 -122 -221 -88
rect -163 -122 -153 -88
rect -91 -122 -85 -88
rect -19 -122 -17 -88
rect 17 -122 19 -88
rect 85 -122 91 -88
rect 153 -122 163 -88
rect 221 -122 235 -88
rect 289 -122 307 -88
rect 357 -122 379 -88
rect 425 -122 451 -88
rect 493 -122 523 -88
rect 561 -122 595 -88
rect 629 -122 663 -88
rect 701 -122 731 -88
rect 773 -122 800 -88
rect 946 -119 980 -85
rect -980 -226 -946 -153
rect 946 -226 980 -153
rect -980 -260 -867 -226
rect -833 -260 -799 -226
rect -765 -260 -731 -226
rect -697 -260 -663 -226
rect -629 -260 -595 -226
rect -561 -260 -527 -226
rect -493 -260 -459 -226
rect -425 -260 -391 -226
rect -357 -260 -323 -226
rect -289 -260 -255 -226
rect -221 -260 -187 -226
rect -153 -260 -119 -226
rect -85 -260 -51 -226
rect -17 -260 17 -226
rect 51 -260 85 -226
rect 119 -260 153 -226
rect 187 -260 221 -226
rect 255 -260 289 -226
rect 323 -260 357 -226
rect 391 -260 425 -226
rect 459 -260 493 -226
rect 527 -260 561 -226
rect 595 -260 629 -226
rect 663 -260 697 -226
rect 731 -260 765 -226
rect 799 -260 833 -226
rect 867 -260 980 -226
<< viali >>
rect -917 226 -883 260
rect -845 226 -833 260
rect -833 226 -811 260
rect -773 226 -765 260
rect -765 226 -739 260
rect -701 226 -697 260
rect -697 226 -667 260
rect -629 226 -595 260
rect -557 226 -527 260
rect -527 226 -523 260
rect -485 226 -459 260
rect -459 226 -451 260
rect -413 226 -391 260
rect -391 226 -379 260
rect -341 226 -323 260
rect -323 226 -307 260
rect -269 226 -255 260
rect -255 226 -235 260
rect -197 226 -187 260
rect -187 226 -163 260
rect -125 226 -119 260
rect -119 226 -91 260
rect -53 226 -51 260
rect -51 226 -19 260
rect 19 226 51 260
rect 51 226 53 260
rect 91 226 119 260
rect 119 226 125 260
rect 163 226 187 260
rect 187 226 197 260
rect 235 226 255 260
rect 255 226 269 260
rect 307 226 323 260
rect 323 226 341 260
rect 379 226 391 260
rect 391 226 413 260
rect 451 226 459 260
rect 459 226 485 260
rect 523 226 527 260
rect 527 226 557 260
rect 595 226 629 260
rect 667 226 697 260
rect 697 226 701 260
rect 739 226 765 260
rect 765 226 773 260
rect 811 226 833 260
rect 833 226 845 260
rect 883 226 917 260
rect -773 88 -765 122
rect -765 88 -739 122
rect -701 88 -697 122
rect -697 88 -667 122
rect -629 88 -595 122
rect -557 88 -527 122
rect -527 88 -523 122
rect -485 88 -459 122
rect -459 88 -451 122
rect -413 88 -391 122
rect -391 88 -379 122
rect -341 88 -323 122
rect -323 88 -307 122
rect -269 88 -255 122
rect -255 88 -235 122
rect -197 88 -187 122
rect -187 88 -163 122
rect -125 88 -119 122
rect -119 88 -91 122
rect -53 88 -51 122
rect -51 88 -19 122
rect 19 88 51 122
rect 51 88 53 122
rect 91 88 119 122
rect 119 88 125 122
rect 163 88 187 122
rect 187 88 197 122
rect 235 88 255 122
rect 255 88 269 122
rect 307 88 323 122
rect 323 88 341 122
rect 379 88 391 122
rect 391 88 413 122
rect 451 88 459 122
rect 459 88 485 122
rect 523 88 527 122
rect 527 88 557 122
rect 595 88 629 122
rect 667 88 697 122
rect 697 88 701 122
rect 739 88 765 122
rect 765 88 773 122
rect -846 -17 -812 17
rect 812 -17 846 17
rect -773 -122 -765 -88
rect -765 -122 -739 -88
rect -701 -122 -697 -88
rect -697 -122 -667 -88
rect -629 -122 -595 -88
rect -557 -122 -527 -88
rect -527 -122 -523 -88
rect -485 -122 -459 -88
rect -459 -122 -451 -88
rect -413 -122 -391 -88
rect -391 -122 -379 -88
rect -341 -122 -323 -88
rect -323 -122 -307 -88
rect -269 -122 -255 -88
rect -255 -122 -235 -88
rect -197 -122 -187 -88
rect -187 -122 -163 -88
rect -125 -122 -119 -88
rect -119 -122 -91 -88
rect -53 -122 -51 -88
rect -51 -122 -19 -88
rect 19 -122 51 -88
rect 51 -122 53 -88
rect 91 -122 119 -88
rect 119 -122 125 -88
rect 163 -122 187 -88
rect 187 -122 197 -88
rect 235 -122 255 -88
rect 255 -122 269 -88
rect 307 -122 323 -88
rect 323 -122 341 -88
rect 379 -122 391 -88
rect 391 -122 413 -88
rect 451 -122 459 -88
rect 459 -122 485 -88
rect 523 -122 527 -88
rect 527 -122 557 -88
rect 595 -122 629 -88
rect 667 -122 697 -88
rect 697 -122 701 -88
rect 739 -122 765 -88
rect 765 -122 773 -88
<< metal1 >>
rect -958 260 958 266
rect -958 226 -917 260
rect -883 226 -845 260
rect -811 226 -773 260
rect -739 226 -701 260
rect -667 226 -629 260
rect -595 226 -557 260
rect -523 226 -485 260
rect -451 226 -413 260
rect -379 226 -341 260
rect -307 226 -269 260
rect -235 226 -197 260
rect -163 226 -125 260
rect -91 226 -53 260
rect -19 226 19 260
rect 53 226 91 260
rect 125 226 163 260
rect 197 226 235 260
rect 269 226 307 260
rect 341 226 379 260
rect 413 226 451 260
rect 485 226 523 260
rect 557 226 595 260
rect 629 226 667 260
rect 701 226 739 260
rect 773 226 811 260
rect 845 226 883 260
rect 917 226 958 260
rect -958 220 958 226
rect -796 122 796 128
rect -796 88 -773 122
rect -739 88 -701 122
rect -667 88 -629 122
rect -595 88 -557 122
rect -523 88 -485 122
rect -451 88 -413 122
rect -379 88 -341 122
rect -307 88 -269 122
rect -235 88 -197 122
rect -163 88 -125 122
rect -91 88 -53 122
rect -19 88 19 122
rect 53 88 91 122
rect 125 88 163 122
rect 197 88 235 122
rect 269 88 307 122
rect 341 88 379 122
rect 413 88 451 122
rect 485 88 523 122
rect 557 88 595 122
rect 629 88 667 122
rect 701 88 739 122
rect 773 88 796 122
rect -796 82 796 88
rect -852 17 -806 50
rect -852 -17 -846 17
rect -812 -17 -806 17
rect -852 -50 -806 -17
rect 806 17 852 50
rect 806 -17 812 17
rect 846 -17 852 17
rect 806 -50 852 -17
rect -796 -88 796 -82
rect -796 -122 -773 -88
rect -739 -122 -701 -88
rect -667 -122 -629 -88
rect -595 -122 -557 -88
rect -523 -122 -485 -88
rect -451 -122 -413 -88
rect -379 -122 -341 -88
rect -307 -122 -269 -88
rect -235 -122 -197 -88
rect -163 -122 -125 -88
rect -91 -122 -53 -88
rect -19 -122 19 -88
rect 53 -122 91 -88
rect 125 -122 163 -88
rect 197 -122 235 -88
rect 269 -122 307 -88
rect 341 -122 379 -88
rect 413 -122 451 -88
rect 485 -122 523 -88
rect 557 -122 595 -88
rect 629 -122 667 -88
rect 701 -122 739 -88
rect 773 -122 796 -88
rect -796 -128 796 -122
<< properties >>
string FIXED_BBOX -963 -243 963 243
<< end >>
