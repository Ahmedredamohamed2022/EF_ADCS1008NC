magic
tech sky130A
magscale 1 2
timestamp 1694078038
<< checkpaint >>
rect -4474 -2252 34066 98074
<< metal1 >>
rect 816 91857 1024 91878
rect 816 91037 859 91857
rect 975 91037 1024 91857
rect 816 91002 1024 91037
rect 4252 91807 4454 91856
rect 4252 91051 4287 91807
rect 4403 91051 4454 91807
rect 7600 91831 7810 91862
rect 14420 91848 14614 91860
rect 7600 91139 7610 91831
rect 7790 91139 7810 91831
rect 7600 91088 7810 91139
rect 11030 91823 11240 91840
rect 11030 91131 11045 91823
rect 11225 91131 11240 91823
rect 14420 91220 14461 91848
rect 14577 91220 14614 91848
rect 17846 91794 18044 91846
rect 17846 91238 17850 91794
rect 14420 91202 14614 91220
rect 18030 91238 18044 91794
rect 21198 91825 21408 91862
rect 17850 91202 18030 91230
rect 11030 91112 11240 91131
rect 21198 91133 21202 91825
rect 21382 91133 21408 91825
rect 21198 91086 21408 91133
rect 24644 91793 24846 91842
rect 24644 91165 24680 91793
rect 24796 91165 24846 91793
rect 24644 91112 24846 91165
rect 4252 91004 4454 91051
rect 816 90988 1018 91002
rect -3018 87645 -1140 87702
rect -3018 87529 -2955 87645
rect -1175 87529 -1140 87645
rect -3018 87434 -1140 87529
rect -628 81992 120 82022
rect -628 81812 -600 81992
rect 92 81812 120 81992
rect -628 81782 120 81812
rect -804 81201 -398 81220
rect -804 81021 -759 81201
rect -451 81021 -398 81201
rect -804 81002 -398 81021
rect -943 78534 -330 78588
rect -943 78516 -226 78534
rect -943 78336 -881 78516
rect -253 78336 -226 78516
rect -943 78318 -226 78336
rect -943 78266 -330 78318
rect -1538 78052 -392 78122
rect -1538 77488 -1476 78052
rect -464 77488 -392 78052
rect -1538 77410 -392 77488
rect -3004 77312 -1532 77330
rect -3004 77132 -2931 77312
rect -1599 77306 -1532 77312
rect -1599 77132 -222 77306
rect -3004 77104 -222 77132
rect -3004 77078 -1532 77104
rect -1044 76956 -268 76980
rect -1046 76938 870 76956
rect -1046 76822 -1022 76938
rect -330 76822 870 76938
rect -1046 76756 870 76822
rect 18712 76839 19260 76886
rect 18712 76723 18771 76839
rect 19207 76723 19260 76839
rect 18712 76682 19260 76723
rect 1172 64248 1284 64656
rect 10330 64559 10432 64592
rect 10330 64507 10353 64559
rect 10405 64507 10432 64559
rect 10330 64495 10432 64507
rect 10330 64443 10353 64495
rect 10405 64443 10432 64495
rect 10330 64431 10432 64443
rect 10330 64404 10353 64431
rect 7864 64379 10353 64404
rect 10405 64379 10432 64431
rect 7864 64367 10432 64379
rect 7864 64315 10353 64367
rect 10405 64315 10432 64367
rect 7864 64303 10432 64315
rect 7864 64251 10353 64303
rect 10405 64251 10432 64303
rect 7864 64239 10432 64251
rect 7864 64187 10353 64239
rect 10405 64187 10432 64239
rect 7864 64184 10432 64187
rect 10330 64175 10432 64184
rect 10330 64123 10353 64175
rect 10405 64123 10432 64175
rect 10330 64111 10432 64123
rect 10330 64059 10353 64111
rect 10405 64059 10432 64111
rect 10330 64026 10432 64059
rect -3144 63574 1282 63608
rect -3144 63458 -3122 63574
rect -2622 63458 1282 63574
rect -3144 63406 1282 63458
rect 28598 63068 31842 63100
rect 28598 62952 31425 63068
rect 31797 62952 31842 63068
rect 28598 62900 31842 62952
rect 10128 57786 10236 57832
rect 10128 57734 10154 57786
rect 10206 57734 10236 57786
rect 10128 57722 10236 57734
rect 10128 57670 10154 57722
rect 10206 57670 10236 57722
rect 7858 57658 10236 57670
rect 7858 57606 10154 57658
rect 10206 57606 10236 57658
rect 7858 57594 10236 57606
rect 7858 57542 10154 57594
rect 10206 57542 10236 57594
rect 7858 57530 10236 57542
rect 7858 57478 10154 57530
rect 10206 57478 10236 57530
rect 7858 57466 10236 57478
rect 7858 57450 10154 57466
rect 10128 57414 10154 57450
rect 10206 57414 10236 57466
rect 10128 57402 10236 57414
rect 10128 57350 10154 57402
rect 10206 57350 10236 57402
rect 10128 57314 10236 57350
rect 1162 56836 1274 57244
rect 17156 57031 17362 57256
rect 10761 56988 18581 57031
rect 10761 56872 10782 56988
rect 11474 56872 18581 56988
rect 10761 56825 18581 56872
rect 23486 56772 23680 57299
rect 26640 56868 26836 57301
rect 26592 56817 27174 56868
rect 23470 56698 23944 56772
rect 23470 56454 23547 56698
rect 23855 56454 23944 56698
rect 26592 56637 26631 56817
rect 27131 56637 27174 56817
rect 26592 56592 27174 56637
rect -3140 56371 1278 56408
rect 23470 56400 23944 56454
rect -3140 56255 -3095 56371
rect -2659 56255 1278 56371
rect -3140 56214 1278 56255
rect 10326 51182 10434 51206
rect 10326 51130 10349 51182
rect 10401 51130 10434 51182
rect 10326 51118 10434 51130
rect 9936 51032 10036 51080
rect 9936 50980 9955 51032
rect 10007 50980 10036 51032
rect 9936 50968 10036 50980
rect 9936 50916 9955 50968
rect 10007 50916 10036 50968
rect 9936 50912 10036 50916
rect 10326 51066 10349 51118
rect 10401 51066 10434 51118
rect 10326 51054 10434 51066
rect 10326 51002 10349 51054
rect 10401 51036 10434 51054
rect 10401 51002 11794 51036
rect 10326 50990 11794 51002
rect 10326 50938 10349 50990
rect 10401 50938 11794 50990
rect 10326 50926 11794 50938
rect 7844 50904 10042 50912
rect 7844 50852 9955 50904
rect 10007 50852 10042 50904
rect 7844 50840 10042 50852
rect 7844 50788 9955 50840
rect 10007 50788 10042 50840
rect 1140 50406 1252 50786
rect 7844 50776 10042 50788
rect 7844 50724 9955 50776
rect 10007 50724 10042 50776
rect 7844 50712 10042 50724
rect 7844 50692 9955 50712
rect 9936 50660 9955 50692
rect 10007 50692 10042 50712
rect 10326 50874 10349 50926
rect 10401 50874 11794 50926
rect 10326 50862 11794 50874
rect 10326 50810 10349 50862
rect 10401 50848 11794 50862
rect 10401 50810 10434 50848
rect 10326 50798 10434 50810
rect 10326 50746 10349 50798
rect 10401 50746 10434 50798
rect 10326 50710 10434 50746
rect 10007 50660 10036 50692
rect 9936 50648 10036 50660
rect 9936 50596 9955 50648
rect 10007 50596 10036 50648
rect 9936 50568 10036 50596
rect -3126 50358 1274 50406
rect -3126 50242 -3097 50358
rect -2661 50242 1274 50358
rect -3126 50196 1274 50242
rect 10126 48406 10232 48466
rect 10126 48354 10154 48406
rect 10206 48354 10232 48406
rect 10126 48342 10232 48354
rect 10126 48290 10154 48342
rect 10206 48290 11772 48342
rect 10126 48278 11772 48290
rect 10126 48226 10154 48278
rect 10206 48226 11772 48278
rect 10126 48214 11772 48226
rect 10126 48162 10154 48214
rect 10206 48162 11772 48214
rect 10126 48150 11772 48162
rect 10126 48098 10154 48150
rect 10206 48126 11772 48150
rect 10206 48098 10232 48126
rect 10126 48086 10232 48098
rect 10126 48034 10154 48086
rect 10206 48034 10232 48086
rect 10126 47994 10232 48034
rect 9512 45752 9620 45792
rect 9512 45700 9540 45752
rect 9592 45700 9620 45752
rect 9512 45688 9620 45700
rect 9512 45636 9540 45688
rect 9592 45636 9620 45688
rect 9512 45624 9620 45636
rect 9512 45572 9540 45624
rect 9592 45614 9620 45624
rect 9592 45572 11460 45614
rect 9512 45560 11460 45572
rect 9512 45508 9540 45560
rect 9592 45508 11460 45560
rect 9512 45496 11460 45508
rect 9512 45444 9540 45496
rect 9592 45458 11460 45496
rect 9592 45444 9620 45458
rect 9512 45432 9620 45444
rect 9512 45380 9540 45432
rect 9592 45380 9620 45432
rect 9512 45342 9620 45380
rect 9730 44276 9836 44314
rect 9730 44224 9756 44276
rect 9808 44224 9836 44276
rect 1126 44016 1238 44218
rect 9730 44212 9836 44224
rect 9730 44160 9756 44212
rect 9808 44160 9836 44212
rect 9730 44148 9836 44160
rect 9730 44142 9756 44148
rect -3110 43991 1238 44016
rect -3110 43811 -3068 43991
rect -2632 43811 1238 43991
rect 7818 44096 9756 44142
rect 9808 44142 9836 44148
rect 9808 44096 9842 44142
rect 7818 44084 9842 44096
rect 7818 44032 9756 44084
rect 9808 44032 9842 44084
rect 7818 44020 9842 44032
rect 7818 43968 9756 44020
rect 9808 43968 9842 44020
rect 7818 43956 9842 43968
rect 7818 43922 9756 43956
rect -3110 43810 1238 43811
rect 9730 43904 9756 43922
rect 9808 43922 9842 43956
rect 9808 43904 9836 43922
rect 9730 43892 9836 43904
rect 9730 43840 9756 43892
rect 9808 43840 9836 43892
rect -3110 43792 1232 43810
rect 9730 43798 9836 43840
rect 9732 42970 9840 43000
rect 9732 42918 9758 42970
rect 9810 42918 9840 42970
rect 9732 42906 9840 42918
rect 9732 42854 9758 42906
rect 9810 42854 9840 42906
rect 9732 42842 9840 42854
rect 9732 42790 9758 42842
rect 9810 42790 9840 42842
rect 9732 42784 9840 42790
rect 9732 42778 11282 42784
rect 9732 42726 9758 42778
rect 9810 42726 11282 42778
rect 9732 42714 11282 42726
rect 9732 42662 9758 42714
rect 9810 42664 11282 42714
rect 9810 42662 9840 42664
rect 9732 42650 9840 42662
rect 9732 42598 9758 42650
rect 9810 42598 9840 42650
rect 9732 42586 9840 42598
rect 9732 42534 9758 42586
rect 9810 42534 9840 42586
rect 9732 42500 9840 42534
rect 9930 40171 10044 40198
rect 9930 40119 9964 40171
rect 10016 40119 10044 40171
rect 9930 40107 10044 40119
rect 9930 40055 9964 40107
rect 10016 40055 10044 40107
rect 9930 40043 10044 40055
rect 9930 40014 9964 40043
rect 9928 39991 9964 40014
rect 10016 40014 10044 40043
rect 10016 39991 11456 40014
rect 9928 39979 11456 39991
rect 9928 39927 9964 39979
rect 10016 39927 11456 39979
rect 9928 39915 11456 39927
rect 9928 39866 9964 39915
rect 9930 39863 9964 39866
rect 10016 39866 11456 39915
rect 10016 39863 10044 39866
rect 9930 39851 10044 39863
rect 9930 39799 9964 39851
rect 10016 39799 10044 39851
rect 9930 39774 10044 39799
rect 9506 37439 9624 37498
rect 9506 37388 9542 37439
rect 7864 37387 9542 37388
rect 9594 37388 9624 37439
rect 9594 37387 9628 37388
rect 7864 37375 9628 37387
rect 7864 37323 9542 37375
rect 9594 37323 9628 37375
rect 7864 37311 9628 37323
rect 7864 37259 9542 37311
rect 9594 37259 9628 37311
rect 7864 37247 9628 37259
rect 7864 37195 9542 37247
rect 9594 37195 9628 37247
rect 7864 37183 9628 37195
rect 1146 37050 1258 37174
rect 7864 37168 9542 37183
rect 9506 37131 9542 37168
rect 9594 37168 9628 37183
rect 9594 37131 9624 37168
rect 9506 37086 9624 37131
rect -3126 37019 1262 37050
rect -3126 36839 -3077 37019
rect -2641 36839 1262 37019
rect -3126 36794 1262 36839
rect 1146 36766 1258 36794
rect 1162 30628 1274 30852
rect -3114 30601 1282 30628
rect -3114 30421 -3092 30601
rect -2592 30421 1282 30601
rect 9312 30555 9426 30594
rect 9312 30503 9338 30555
rect 9390 30503 9426 30555
rect 9312 30491 9426 30503
rect 9312 30446 9338 30491
rect -3114 30380 1282 30421
rect 7868 30439 9338 30446
rect 9390 30439 9426 30491
rect 7868 30427 9426 30439
rect 7868 30375 9338 30427
rect 9390 30375 9426 30427
rect 7868 30363 9426 30375
rect 7868 30311 9338 30363
rect 9390 30311 9426 30363
rect 7868 30299 9426 30311
rect 7868 30247 9338 30299
rect 9390 30247 9426 30299
rect 7868 30235 9426 30247
rect 7868 30226 9338 30235
rect 9312 30183 9338 30226
rect 9390 30183 9426 30235
rect 9312 30136 9426 30183
rect 9310 25977 9418 26020
rect 9310 25925 9338 25977
rect 9390 25925 9418 25977
rect 9310 25913 9418 25925
rect 9310 25861 9338 25913
rect 9390 25861 9418 25913
rect 9310 25849 9418 25861
rect 9310 25797 9338 25849
rect 9390 25840 9418 25849
rect 9390 25797 11452 25840
rect 9310 25785 11452 25797
rect 9310 25733 9338 25785
rect 9390 25733 11452 25785
rect 9310 25721 11452 25733
rect 9310 25669 9338 25721
rect 9390 25669 11452 25721
rect 9310 25657 11452 25669
rect 9310 25605 9338 25657
rect 9390 25652 11452 25657
rect 9390 25605 9418 25652
rect 9310 25560 9418 25605
rect 1140 23820 1252 23878
rect -3104 23772 1252 23820
rect -3104 23656 -3030 23772
rect -2658 23656 1252 23772
rect 9078 23821 9224 23852
rect 9078 23769 9114 23821
rect 9166 23769 9224 23821
rect 9078 23757 9224 23769
rect 9078 23705 9114 23757
rect 9166 23705 9224 23757
rect 9078 23702 9224 23705
rect -3104 23584 1252 23656
rect 1140 23470 1252 23584
rect 7854 23693 9224 23702
rect 7854 23641 9114 23693
rect 9166 23641 9224 23693
rect 7854 23629 9224 23641
rect 7854 23577 9114 23629
rect 9166 23577 9224 23629
rect 7854 23565 9224 23577
rect 7854 23513 9114 23565
rect 9166 23513 9224 23565
rect 7854 23501 9224 23513
rect 7854 23482 9114 23501
rect 9078 23449 9114 23482
rect 9166 23449 9224 23501
rect 9078 23146 9224 23449
rect 9078 22936 11524 23146
rect 9088 22930 11524 22936
rect 8488 20650 8644 20694
rect 8488 20598 8517 20650
rect 8569 20598 8644 20650
rect 8488 20586 8644 20598
rect 8488 20534 8517 20586
rect 8569 20534 8644 20586
rect 8488 20522 8644 20534
rect 8488 20470 8517 20522
rect 8569 20470 8644 20522
rect 8488 20458 8644 20470
rect 8488 20406 8517 20458
rect 8569 20418 8644 20458
rect 8569 20406 11492 20418
rect 8488 20394 11492 20406
rect 8488 20342 8517 20394
rect 8569 20342 11492 20394
rect 8488 20330 11492 20342
rect 8488 20278 8517 20330
rect 8569 20278 11492 20330
rect 8488 20266 11492 20278
rect 8488 20214 8517 20266
rect 8569 20262 11492 20266
rect 8569 20214 8644 20262
rect 8488 20202 8644 20214
rect 8488 20150 8517 20202
rect 8569 20150 8644 20202
rect 8488 20138 8644 20150
rect 8488 20086 8517 20138
rect 8569 20086 8644 20138
rect 8488 20074 8644 20086
rect 8488 20022 8517 20074
rect 8569 20022 8644 20074
rect 8488 19984 8644 20022
rect 8702 17748 8822 17802
rect 8702 17696 8727 17748
rect 8779 17696 8822 17748
rect 8702 17684 8822 17696
rect 8702 17632 8727 17684
rect 8779 17632 8822 17684
rect 8702 17620 8822 17632
rect 8702 17568 8727 17620
rect 8779 17588 8822 17620
rect 8779 17568 11518 17588
rect 8702 17556 11518 17568
rect 8702 17504 8727 17556
rect 8779 17504 11518 17556
rect 8702 17492 11518 17504
rect 8702 17440 8727 17492
rect 8779 17468 11518 17492
rect 8779 17440 8822 17468
rect 8702 17428 8822 17440
rect 8702 17376 8727 17428
rect 8779 17376 8822 17428
rect 8702 17364 8822 17376
rect 8702 17312 8727 17364
rect 8779 17312 8822 17364
rect 8702 17300 8822 17312
rect 8702 17248 8727 17300
rect 8779 17248 8822 17300
rect 8702 17198 8822 17248
rect 8906 17001 9002 17036
rect 8906 16949 8932 17001
rect 8984 16949 9002 17001
rect 8906 16937 9002 16949
rect 1146 16812 1258 16926
rect 8906 16896 8932 16937
rect -3100 16768 1258 16812
rect -3100 16652 -3046 16768
rect -2674 16652 1258 16768
rect 7854 16885 8932 16896
rect 8984 16896 9002 16937
rect 8984 16885 9008 16896
rect 7854 16873 9008 16885
rect 7854 16821 8932 16873
rect 8984 16821 9008 16873
rect 7854 16809 9008 16821
rect 7854 16757 8932 16809
rect 8984 16757 9008 16809
rect 7854 16745 9008 16757
rect 7854 16693 8932 16745
rect 8984 16693 9008 16745
rect 7854 16681 9008 16693
rect 7854 16676 8932 16681
rect -3100 16594 1258 16652
rect 8906 16629 8932 16676
rect 8984 16676 9008 16681
rect 8984 16629 9002 16676
rect 8906 16600 9002 16629
rect 1146 16518 1258 16594
rect 8904 14969 9052 15024
rect 8904 14917 8927 14969
rect 8979 14917 9052 14969
rect 8904 14905 9052 14917
rect 8904 14853 8927 14905
rect 8979 14853 9052 14905
rect 8904 14841 9052 14853
rect 8904 14789 8927 14841
rect 8979 14818 9052 14841
rect 8979 14789 11384 14818
rect 8904 14777 11384 14789
rect 8904 14725 8927 14777
rect 8979 14725 11384 14777
rect 8904 14713 11384 14725
rect 8904 14661 8927 14713
rect 8979 14670 11384 14713
rect 8979 14661 9052 14670
rect 8904 14649 9052 14661
rect 8904 14597 8927 14649
rect 8979 14597 9052 14649
rect 8904 14585 9052 14597
rect 8904 14533 8927 14585
rect 8979 14533 9052 14585
rect 8904 14488 9052 14533
rect 8698 10437 8804 10526
rect 8698 10385 8722 10437
rect 8774 10385 8804 10437
rect 8698 10373 8804 10385
rect 8698 10342 8722 10373
rect 7834 10321 8722 10342
rect 8774 10342 8804 10373
rect 8774 10321 8808 10342
rect 7834 10309 8808 10321
rect 7834 10257 8722 10309
rect 8774 10257 8808 10309
rect 7834 10245 8808 10257
rect 7834 10193 8722 10245
rect 8774 10193 8808 10245
rect 7834 10181 8808 10193
rect 7834 10129 8722 10181
rect 8774 10129 8808 10181
rect 7834 10122 8808 10129
rect 8698 10117 8804 10122
rect 8698 10065 8722 10117
rect 8774 10065 8804 10117
rect 8698 10022 8804 10065
rect -3092 9978 1239 10020
rect -3092 9862 -3052 9978
rect -2552 9862 1239 9978
rect -3092 9798 1239 9862
rect 7854 3339 8592 3388
rect 7854 3223 8419 3339
rect 8535 3223 8592 3339
rect 7854 3168 8592 3223
rect -3050 2773 1260 2814
rect -3050 2657 -2994 2773
rect -2558 2657 1260 2773
rect -3050 2590 1260 2657
rect 1620 1346 2088 1394
rect 1620 1102 1663 1346
rect 2035 1102 2088 1346
rect 1620 1018 2088 1102
<< via1 >>
rect 859 91037 975 91857
rect 4287 91051 4403 91807
rect 7610 91139 7790 91831
rect 11045 91131 11225 91823
rect 14461 91220 14577 91848
rect 17850 91230 18030 91794
rect 21202 91133 21382 91825
rect 24680 91165 24796 91793
rect -2955 87529 -1175 87645
rect -600 81812 92 81992
rect -759 81021 -451 81201
rect -881 78336 -253 78516
rect -1476 77488 -464 78052
rect -2931 77132 -1599 77312
rect -1022 76822 -330 76938
rect 18771 76723 19207 76839
rect 10353 64507 10405 64559
rect 10353 64443 10405 64495
rect 10353 64379 10405 64431
rect 10353 64315 10405 64367
rect 10353 64251 10405 64303
rect 10353 64187 10405 64239
rect 10353 64123 10405 64175
rect 10353 64059 10405 64111
rect -3122 63458 -2622 63574
rect 31425 62952 31797 63068
rect 10154 57734 10206 57786
rect 10154 57670 10206 57722
rect 10154 57606 10206 57658
rect 10154 57542 10206 57594
rect 10154 57478 10206 57530
rect 10154 57414 10206 57466
rect 10154 57350 10206 57402
rect 10782 56872 11474 56988
rect 23547 56454 23855 56698
rect 26631 56637 27131 56817
rect -3095 56255 -2659 56371
rect 10349 51130 10401 51182
rect 9955 50980 10007 51032
rect 9955 50916 10007 50968
rect 10349 51066 10401 51118
rect 10349 51002 10401 51054
rect 10349 50938 10401 50990
rect 9955 50852 10007 50904
rect 9955 50788 10007 50840
rect 9955 50724 10007 50776
rect 9955 50660 10007 50712
rect 10349 50874 10401 50926
rect 10349 50810 10401 50862
rect 10349 50746 10401 50798
rect 9955 50596 10007 50648
rect -3097 50242 -2661 50358
rect 10154 48354 10206 48406
rect 10154 48290 10206 48342
rect 10154 48226 10206 48278
rect 10154 48162 10206 48214
rect 10154 48098 10206 48150
rect 10154 48034 10206 48086
rect 9540 45700 9592 45752
rect 9540 45636 9592 45688
rect 9540 45572 9592 45624
rect 9540 45508 9592 45560
rect 9540 45444 9592 45496
rect 9540 45380 9592 45432
rect 9756 44224 9808 44276
rect 9756 44160 9808 44212
rect -3068 43811 -2632 43991
rect 9756 44096 9808 44148
rect 9756 44032 9808 44084
rect 9756 43968 9808 44020
rect 9756 43904 9808 43956
rect 9756 43840 9808 43892
rect 9758 42918 9810 42970
rect 9758 42854 9810 42906
rect 9758 42790 9810 42842
rect 9758 42726 9810 42778
rect 9758 42662 9810 42714
rect 9758 42598 9810 42650
rect 9758 42534 9810 42586
rect 9964 40119 10016 40171
rect 9964 40055 10016 40107
rect 9964 39991 10016 40043
rect 9964 39927 10016 39979
rect 9964 39863 10016 39915
rect 9964 39799 10016 39851
rect 9542 37387 9594 37439
rect 9542 37323 9594 37375
rect 9542 37259 9594 37311
rect 9542 37195 9594 37247
rect 9542 37131 9594 37183
rect -3077 36839 -2641 37019
rect -3092 30421 -2592 30601
rect 9338 30503 9390 30555
rect 9338 30439 9390 30491
rect 9338 30375 9390 30427
rect 9338 30311 9390 30363
rect 9338 30247 9390 30299
rect 9338 30183 9390 30235
rect 9338 25925 9390 25977
rect 9338 25861 9390 25913
rect 9338 25797 9390 25849
rect 9338 25733 9390 25785
rect 9338 25669 9390 25721
rect 9338 25605 9390 25657
rect -3030 23656 -2658 23772
rect 9114 23769 9166 23821
rect 9114 23705 9166 23757
rect 9114 23641 9166 23693
rect 9114 23577 9166 23629
rect 9114 23513 9166 23565
rect 9114 23449 9166 23501
rect 8517 20598 8569 20650
rect 8517 20534 8569 20586
rect 8517 20470 8569 20522
rect 8517 20406 8569 20458
rect 8517 20342 8569 20394
rect 8517 20278 8569 20330
rect 8517 20214 8569 20266
rect 8517 20150 8569 20202
rect 8517 20086 8569 20138
rect 8517 20022 8569 20074
rect 8727 17696 8779 17748
rect 8727 17632 8779 17684
rect 8727 17568 8779 17620
rect 8727 17504 8779 17556
rect 8727 17440 8779 17492
rect 8727 17376 8779 17428
rect 8727 17312 8779 17364
rect 8727 17248 8779 17300
rect 8932 16949 8984 17001
rect -3046 16652 -2674 16768
rect 8932 16885 8984 16937
rect 8932 16821 8984 16873
rect 8932 16757 8984 16809
rect 8932 16693 8984 16745
rect 8932 16629 8984 16681
rect 8927 14917 8979 14969
rect 8927 14853 8979 14905
rect 8927 14789 8979 14841
rect 8927 14725 8979 14777
rect 8927 14661 8979 14713
rect 8927 14597 8979 14649
rect 8927 14533 8979 14585
rect 8722 10385 8774 10437
rect 8722 10321 8774 10373
rect 8722 10257 8774 10309
rect 8722 10193 8774 10245
rect 8722 10129 8774 10181
rect 8722 10065 8774 10117
rect -3052 9862 -2552 9978
rect 8419 3223 8535 3339
rect -2994 2657 -2558 2773
rect 1663 1102 2035 1346
<< metal2 >>
rect 1152 96524 1346 96802
rect 1152 95998 1351 96524
rect 4582 96516 4794 96806
rect 7924 96560 8136 96806
rect 816 91857 1024 91878
rect 816 91037 859 91857
rect 975 91526 1024 91857
rect 1157 91526 1351 95998
rect 975 91332 1351 91526
rect 4238 91807 4444 91852
rect 975 91037 1024 91332
rect 816 91002 1024 91037
rect 4238 91051 4287 91807
rect 4403 91608 4444 91807
rect 4579 91608 4809 96516
rect 4403 91378 4809 91608
rect 7604 91831 7810 91874
rect 7604 91584 7610 91831
rect 4403 91051 4444 91378
rect 7602 91360 7610 91584
rect 7604 91139 7610 91360
rect 7790 91584 7810 91831
rect 7922 91584 8146 96560
rect 11350 96516 11562 96800
rect 11345 95812 11562 96516
rect 14700 96546 14912 96806
rect 14700 95818 14915 96546
rect 18178 96494 18390 96814
rect 7790 91360 8146 91584
rect 11022 91823 11240 91856
rect 7790 91139 7810 91360
rect 7604 91084 7810 91139
rect 11022 91131 11045 91823
rect 11225 91602 11240 91823
rect 11345 91602 11559 95812
rect 11225 91388 11559 91602
rect 14414 91848 14620 91880
rect 11225 91131 11240 91388
rect 14414 91220 14461 91848
rect 14577 91616 14620 91848
rect 14713 91616 14915 95818
rect 17836 91794 18034 91840
rect 17836 91656 17850 91794
rect 14577 91414 14915 91616
rect 17832 91432 17850 91656
rect 14577 91220 14620 91414
rect 14414 91190 14620 91220
rect 17836 91230 17850 91432
rect 18030 91656 18034 91794
rect 18176 91656 18400 96494
rect 21494 95818 21706 96806
rect 24870 96568 25082 96806
rect 24870 95818 25094 96568
rect 18030 91432 18400 91656
rect 21190 91825 21396 91880
rect 21190 91532 21202 91825
rect 18030 91230 18034 91432
rect 21184 91340 21202 91532
rect 17836 91172 18034 91230
rect 11022 91090 11240 91131
rect 21190 91133 21202 91340
rect 21382 91532 21396 91825
rect 21494 91532 21686 95818
rect 21382 91340 21686 91532
rect 24638 91793 24844 91844
rect 21382 91133 21396 91340
rect 21190 91094 21396 91133
rect 24638 91165 24680 91793
rect 24796 91564 24844 91793
rect 24878 91564 25094 95818
rect 24796 91348 25094 91564
rect 24796 91165 24844 91348
rect 24638 91124 24844 91165
rect 4238 91010 4444 91051
rect -3020 87655 -1118 87692
rect -3020 87645 -2933 87655
rect -1197 87645 -1118 87655
rect -3020 87529 -2955 87645
rect -1175 87529 -1118 87645
rect -3020 87519 -2933 87529
rect -1197 87519 -1118 87529
rect -3020 87440 -1118 87519
rect -2070 86506 -1638 86542
rect -2070 86130 -2005 86506
rect -1709 86130 -1638 86506
rect -2070 78122 -1638 86130
rect -1470 85885 -1174 85928
rect -1470 85509 -1434 85885
rect -1218 85509 -1174 85885
rect -1470 78584 -1174 85509
rect 25156 85863 25632 91680
rect 25156 85567 25223 85863
rect 25599 85567 25632 85863
rect 25156 85488 25632 85567
rect 29790 85846 30422 85924
rect 29790 85550 29832 85846
rect 30368 85550 30422 85846
rect -1064 85137 -748 85210
rect -1064 84841 -1019 85137
rect -803 84841 -748 85137
rect -1064 82066 -748 84841
rect 24826 85165 25331 85212
rect 24826 84789 24852 85165
rect 25308 84789 25331 85165
rect 24826 83768 25331 84789
rect 25726 84571 26404 84638
rect 25726 84435 25761 84571
rect 26377 84435 26404 84571
rect 25726 84374 26404 84435
rect 26009 83627 26088 84374
rect 29790 83584 30422 85550
rect -658 82066 174 82070
rect -1064 81992 174 82066
rect -1064 81812 -600 81992
rect 92 81812 174 81992
rect -1064 81750 174 81812
rect -658 81740 174 81750
rect -804 81201 -398 81220
rect -804 81021 -759 81201
rect -451 81021 -398 81201
rect -804 81002 -398 81021
rect -944 78584 -186 78590
rect -1470 78516 -186 78584
rect -1470 78336 -881 78516
rect -253 78336 -186 78516
rect -1470 78282 -186 78336
rect -944 78278 -186 78282
rect -2070 78052 -392 78122
rect -2070 77488 -1476 78052
rect -464 77488 -392 78052
rect -2070 77412 -392 77488
rect -1770 77410 -392 77412
rect -3004 77114 -2933 77330
rect -1597 77114 -1532 77330
rect -3004 77078 -1532 77114
rect -1044 76948 -268 76980
rect -1044 76812 -1024 76948
rect -328 76812 -268 76948
rect 19100 76886 19320 76888
rect -1044 76756 -268 76812
rect 18712 76839 19320 76886
rect 18712 76786 18771 76839
rect 18710 76723 18771 76786
rect 19207 76723 19320 76839
rect 18710 76686 19320 76723
rect 18712 76682 19320 76686
rect 19100 72160 19320 76682
rect 26980 72160 27200 72792
rect 19100 71940 27200 72160
rect 27246 71740 27466 72714
rect 26836 71736 26898 71740
rect 27208 71736 27470 71740
rect 17228 71516 27470 71736
rect -3138 63584 -2588 63616
rect -3138 63574 -3100 63584
rect -2644 63574 -2588 63584
rect -3138 63458 -3122 63574
rect -2622 63458 -2588 63574
rect -3138 63448 -3100 63458
rect -2644 63448 -2588 63458
rect -3138 63406 -2588 63448
rect -3144 56381 -2598 56408
rect -3144 56245 -3105 56381
rect -2649 56245 -2598 56381
rect -3144 56210 -2598 56245
rect -3134 50368 -2588 50394
rect -3134 50232 -3107 50368
rect -2651 50232 -2588 50368
rect -3134 50188 -2588 50232
rect -3114 43991 -2584 44020
rect -3114 43969 -3068 43991
rect -2632 43969 -2584 43991
rect -3114 43833 -3078 43969
rect -2622 43833 -2584 43969
rect -3114 43811 -3068 43833
rect -2632 43811 -2584 43833
rect -3114 43788 -2584 43811
rect -3122 37019 -2584 37046
rect -3122 36839 -3077 37019
rect -2641 36839 -2584 37019
rect -3122 36794 -2584 36839
rect -3122 30619 -2562 30634
rect -3122 30601 -3070 30619
rect -2614 30601 -2562 30619
rect -3122 30421 -3092 30601
rect -2592 30421 -2562 30601
rect -3122 30403 -3070 30421
rect -2614 30403 -2562 30421
rect -3122 30384 -2562 30403
rect -3100 23782 -2596 23824
rect -3100 23646 -3032 23782
rect -2656 23646 -2596 23782
rect -3100 23604 -2596 23646
rect 8498 20650 8602 65646
rect 8498 20598 8517 20650
rect 8569 20598 8602 20650
rect 8498 20586 8602 20598
rect 8498 20534 8517 20586
rect 8569 20534 8602 20586
rect 8498 20522 8602 20534
rect 8498 20470 8517 20522
rect 8569 20470 8602 20522
rect 8498 20458 8602 20470
rect 8498 20406 8517 20458
rect 8569 20406 8602 20458
rect 8498 20394 8602 20406
rect 8498 20342 8517 20394
rect 8569 20342 8602 20394
rect 8498 20330 8602 20342
rect 8498 20278 8517 20330
rect 8569 20278 8602 20330
rect 8498 20266 8602 20278
rect 8498 20214 8517 20266
rect 8569 20214 8602 20266
rect 8498 20202 8602 20214
rect 8498 20150 8517 20202
rect 8569 20150 8602 20202
rect 8498 20138 8602 20150
rect 8498 20086 8517 20138
rect 8569 20086 8602 20138
rect 8498 20074 8602 20086
rect 8498 20022 8517 20074
rect 8569 20022 8602 20074
rect -3096 16778 -2592 16812
rect -3096 16642 -3048 16778
rect -2672 16642 -2592 16778
rect -3096 16602 -2592 16642
rect -3082 9988 -2512 10016
rect -3082 9978 -3030 9988
rect -2574 9978 -2512 9988
rect -3082 9862 -3052 9978
rect -2552 9862 -2512 9978
rect -3082 9852 -3030 9862
rect -2574 9852 -2512 9862
rect -3082 9806 -2512 9852
rect 8498 3388 8602 20022
rect 8372 3339 8602 3388
rect 8372 3223 8419 3339
rect 8535 3223 8602 3339
rect 8372 3168 8602 3223
rect -3054 2783 -2480 2816
rect -3054 2647 -3004 2783
rect -2548 2647 -2480 2783
rect -3054 2598 -2480 2647
rect 1620 1346 2088 1394
rect 1620 1332 1663 1346
rect 2035 1332 2088 1346
rect 1620 1116 1661 1332
rect 2037 1116 2088 1332
rect 1620 1102 1663 1116
rect 2035 1102 2088 1116
rect 1620 1018 2088 1102
rect 8498 652 8602 3168
rect 8700 17748 8804 65646
rect 8700 17696 8727 17748
rect 8779 17696 8804 17748
rect 8700 17684 8804 17696
rect 8700 17632 8727 17684
rect 8779 17632 8804 17684
rect 8700 17620 8804 17632
rect 8700 17568 8727 17620
rect 8779 17568 8804 17620
rect 8700 17556 8804 17568
rect 8700 17504 8727 17556
rect 8779 17504 8804 17556
rect 8700 17492 8804 17504
rect 8700 17440 8727 17492
rect 8779 17440 8804 17492
rect 8700 17428 8804 17440
rect 8700 17376 8727 17428
rect 8779 17376 8804 17428
rect 8700 17364 8804 17376
rect 8700 17312 8727 17364
rect 8779 17312 8804 17364
rect 8700 17300 8804 17312
rect 8700 17248 8727 17300
rect 8779 17248 8804 17300
rect 8700 10437 8804 17248
rect 8700 10385 8722 10437
rect 8774 10385 8804 10437
rect 8700 10373 8804 10385
rect 8700 10321 8722 10373
rect 8774 10321 8804 10373
rect 8700 10309 8804 10321
rect 8700 10257 8722 10309
rect 8774 10257 8804 10309
rect 8700 10245 8804 10257
rect 8700 10193 8722 10245
rect 8774 10193 8804 10245
rect 8700 10181 8804 10193
rect 8700 10129 8722 10181
rect 8774 10129 8804 10181
rect 8700 10117 8804 10129
rect 8700 10065 8722 10117
rect 8774 10065 8804 10117
rect 8700 602 8804 10065
rect 8904 17001 9008 65646
rect 8904 16949 8932 17001
rect 8984 16949 9008 17001
rect 8904 16937 9008 16949
rect 8904 16885 8932 16937
rect 8984 16885 9008 16937
rect 8904 16873 9008 16885
rect 8904 16821 8932 16873
rect 8984 16821 9008 16873
rect 8904 16809 9008 16821
rect 8904 16757 8932 16809
rect 8984 16757 9008 16809
rect 8904 16745 9008 16757
rect 8904 16693 8932 16745
rect 8984 16693 9008 16745
rect 8904 16681 9008 16693
rect 8904 16629 8932 16681
rect 8984 16629 9008 16681
rect 8904 14969 9008 16629
rect 8904 14917 8927 14969
rect 8979 14917 9008 14969
rect 8904 14905 9008 14917
rect 8904 14853 8927 14905
rect 8979 14853 9008 14905
rect 8904 14841 9008 14853
rect 8904 14789 8927 14841
rect 8979 14789 9008 14841
rect 8904 14777 9008 14789
rect 8904 14725 8927 14777
rect 8979 14725 9008 14777
rect 8904 14713 9008 14725
rect 8904 14661 8927 14713
rect 8979 14661 9008 14713
rect 8904 14649 9008 14661
rect 8904 14597 8927 14649
rect 8979 14597 9008 14649
rect 8904 14585 9008 14597
rect 8904 14533 8927 14585
rect 8979 14533 9008 14585
rect 8904 602 9008 14533
rect 9094 23821 9198 65646
rect 9094 23769 9114 23821
rect 9166 23769 9198 23821
rect 9094 23757 9198 23769
rect 9094 23705 9114 23757
rect 9166 23705 9198 23757
rect 9094 23693 9198 23705
rect 9094 23641 9114 23693
rect 9166 23641 9198 23693
rect 9094 23629 9198 23641
rect 9094 23577 9114 23629
rect 9166 23577 9198 23629
rect 9094 23565 9198 23577
rect 9094 23513 9114 23565
rect 9166 23513 9198 23565
rect 9094 23501 9198 23513
rect 9094 23449 9114 23501
rect 9166 23449 9198 23501
rect 9094 602 9198 23449
rect 9316 30555 9420 65646
rect 9316 30503 9338 30555
rect 9390 30503 9420 30555
rect 9316 30491 9420 30503
rect 9316 30439 9338 30491
rect 9390 30439 9420 30491
rect 9316 30427 9420 30439
rect 9316 30375 9338 30427
rect 9390 30375 9420 30427
rect 9316 30363 9420 30375
rect 9316 30311 9338 30363
rect 9390 30311 9420 30363
rect 9316 30299 9420 30311
rect 9316 30247 9338 30299
rect 9390 30247 9420 30299
rect 9316 30235 9420 30247
rect 9316 30183 9338 30235
rect 9390 30183 9420 30235
rect 9316 25977 9420 30183
rect 9316 25925 9338 25977
rect 9390 25925 9420 25977
rect 9316 25913 9420 25925
rect 9316 25861 9338 25913
rect 9390 25861 9420 25913
rect 9316 25849 9420 25861
rect 9316 25797 9338 25849
rect 9390 25797 9420 25849
rect 9316 25785 9420 25797
rect 9316 25733 9338 25785
rect 9390 25733 9420 25785
rect 9316 25721 9420 25733
rect 9316 25669 9338 25721
rect 9390 25669 9420 25721
rect 9316 25657 9420 25669
rect 9316 25605 9338 25657
rect 9390 25605 9420 25657
rect 9316 602 9420 25605
rect 9516 45752 9620 65646
rect 9516 45700 9540 45752
rect 9592 45700 9620 45752
rect 9516 45688 9620 45700
rect 9516 45636 9540 45688
rect 9592 45636 9620 45688
rect 9516 45624 9620 45636
rect 9516 45572 9540 45624
rect 9592 45572 9620 45624
rect 9516 45560 9620 45572
rect 9516 45508 9540 45560
rect 9592 45508 9620 45560
rect 9516 45496 9620 45508
rect 9516 45444 9540 45496
rect 9592 45444 9620 45496
rect 9516 45432 9620 45444
rect 9516 45380 9540 45432
rect 9592 45380 9620 45432
rect 9516 37439 9620 45380
rect 9516 37387 9542 37439
rect 9594 37387 9620 37439
rect 9516 37375 9620 37387
rect 9516 37323 9542 37375
rect 9594 37323 9620 37375
rect 9516 37311 9620 37323
rect 9516 37259 9542 37311
rect 9594 37259 9620 37311
rect 9516 37247 9620 37259
rect 9516 37195 9542 37247
rect 9594 37195 9620 37247
rect 9516 37183 9620 37195
rect 9516 37131 9542 37183
rect 9594 37131 9620 37183
rect 9516 602 9620 37131
rect 9738 44276 9842 65646
rect 9738 44224 9756 44276
rect 9808 44224 9842 44276
rect 9738 44212 9842 44224
rect 9738 44160 9756 44212
rect 9808 44160 9842 44212
rect 9738 44148 9842 44160
rect 9738 44096 9756 44148
rect 9808 44096 9842 44148
rect 9738 44084 9842 44096
rect 9738 44032 9756 44084
rect 9808 44032 9842 44084
rect 9738 44020 9842 44032
rect 9738 43968 9756 44020
rect 9808 43968 9842 44020
rect 9738 43956 9842 43968
rect 9738 43904 9756 43956
rect 9808 43904 9842 43956
rect 9738 43892 9842 43904
rect 9738 43840 9756 43892
rect 9808 43840 9842 43892
rect 9738 42970 9842 43840
rect 9738 42918 9758 42970
rect 9810 42918 9842 42970
rect 9738 42906 9842 42918
rect 9738 42854 9758 42906
rect 9810 42854 9842 42906
rect 9738 42842 9842 42854
rect 9738 42790 9758 42842
rect 9810 42790 9842 42842
rect 9738 42778 9842 42790
rect 9738 42726 9758 42778
rect 9810 42726 9842 42778
rect 9738 42714 9842 42726
rect 9738 42662 9758 42714
rect 9810 42662 9842 42714
rect 9738 42650 9842 42662
rect 9738 42598 9758 42650
rect 9810 42598 9842 42650
rect 9738 42586 9842 42598
rect 9738 42534 9758 42586
rect 9810 42534 9842 42586
rect 9738 602 9842 42534
rect 9936 51032 10040 65646
rect 9936 50980 9955 51032
rect 10007 50980 10040 51032
rect 9936 50968 10040 50980
rect 9936 50916 9955 50968
rect 10007 50916 10040 50968
rect 9936 50904 10040 50916
rect 9936 50852 9955 50904
rect 10007 50852 10040 50904
rect 9936 50840 10040 50852
rect 9936 50788 9955 50840
rect 10007 50788 10040 50840
rect 9936 50776 10040 50788
rect 9936 50724 9955 50776
rect 10007 50724 10040 50776
rect 9936 50712 10040 50724
rect 9936 50660 9955 50712
rect 10007 50660 10040 50712
rect 9936 50648 10040 50660
rect 9936 50596 9955 50648
rect 10007 50596 10040 50648
rect 9936 40171 10040 50596
rect 9936 40119 9964 40171
rect 10016 40119 10040 40171
rect 9936 40107 10040 40119
rect 9936 40055 9964 40107
rect 10016 40055 10040 40107
rect 9936 40043 10040 40055
rect 9936 39991 9964 40043
rect 10016 39991 10040 40043
rect 9936 39979 10040 39991
rect 9936 39927 9964 39979
rect 10016 39927 10040 39979
rect 9936 39915 10040 39927
rect 9936 39863 9964 39915
rect 10016 39863 10040 39915
rect 9936 39851 10040 39863
rect 9936 39799 9964 39851
rect 10016 39799 10040 39851
rect 9936 602 10040 39799
rect 10128 57786 10232 65646
rect 10128 57734 10154 57786
rect 10206 57734 10232 57786
rect 10128 57722 10232 57734
rect 10128 57670 10154 57722
rect 10206 57670 10232 57722
rect 10128 57658 10232 57670
rect 10128 57606 10154 57658
rect 10206 57606 10232 57658
rect 10128 57594 10232 57606
rect 10128 57542 10154 57594
rect 10206 57542 10232 57594
rect 10128 57530 10232 57542
rect 10128 57478 10154 57530
rect 10206 57478 10232 57530
rect 10128 57466 10232 57478
rect 10128 57414 10154 57466
rect 10206 57414 10232 57466
rect 10128 57402 10232 57414
rect 10128 57350 10154 57402
rect 10206 57350 10232 57402
rect 10128 48406 10232 57350
rect 10128 48354 10154 48406
rect 10206 48354 10232 48406
rect 10128 48342 10232 48354
rect 10128 48290 10154 48342
rect 10206 48290 10232 48342
rect 10128 48278 10232 48290
rect 10128 48226 10154 48278
rect 10206 48226 10232 48278
rect 10128 48214 10232 48226
rect 10128 48162 10154 48214
rect 10206 48162 10232 48214
rect 10128 48150 10232 48162
rect 10128 48098 10154 48150
rect 10206 48098 10232 48150
rect 10128 48086 10232 48098
rect 10128 48034 10154 48086
rect 10206 48034 10232 48086
rect 10128 602 10232 48034
rect 10330 64559 10434 65646
rect 10330 64507 10353 64559
rect 10405 64507 10434 64559
rect 10330 64495 10434 64507
rect 10330 64443 10353 64495
rect 10405 64443 10434 64495
rect 10330 64431 10434 64443
rect 10330 64379 10353 64431
rect 10405 64379 10434 64431
rect 10330 64367 10434 64379
rect 10330 64315 10353 64367
rect 10405 64315 10434 64367
rect 10330 64303 10434 64315
rect 10330 64251 10353 64303
rect 10405 64251 10434 64303
rect 10330 64239 10434 64251
rect 10330 64187 10353 64239
rect 10405 64187 10434 64239
rect 10330 64175 10434 64187
rect 10330 64123 10353 64175
rect 10405 64123 10434 64175
rect 10330 64111 10434 64123
rect 10330 64059 10353 64111
rect 10405 64059 10434 64111
rect 10330 51182 10434 64059
rect 17228 64018 17448 71516
rect 31392 63078 31842 63104
rect 31392 62942 31423 63078
rect 31799 62942 31842 63078
rect 31392 62908 31842 62942
rect 15380 57365 16564 57404
rect 15380 57229 15411 57365
rect 16507 57229 16564 57365
rect 15380 57188 16564 57229
rect 10766 56998 11504 57022
rect 10766 56862 10780 56998
rect 11476 56862 11504 56998
rect 10766 56822 11504 56862
rect 16816 56712 17018 57454
rect 17616 57316 18796 57320
rect 17616 57180 17618 57316
rect 18794 57180 18796 57316
rect 17616 57176 18796 57180
rect 26592 56817 27174 56868
rect 16618 56687 17240 56712
rect 16618 56471 16663 56687
rect 17199 56471 17240 56687
rect 16618 56438 17240 56471
rect 23470 56698 23944 56772
rect 23470 56454 23547 56698
rect 23855 56454 23944 56698
rect 26592 56637 26631 56817
rect 27131 56637 27174 56817
rect 26592 56592 27174 56637
rect 23470 56400 23944 56454
rect 10330 51130 10349 51182
rect 10401 51130 10434 51182
rect 10330 51118 10434 51130
rect 10330 51066 10349 51118
rect 10401 51066 10434 51118
rect 10330 51054 10434 51066
rect 10330 51002 10349 51054
rect 10401 51002 10434 51054
rect 10330 50990 10434 51002
rect 10330 50938 10349 50990
rect 10401 50938 10434 50990
rect 10330 50926 10434 50938
rect 10330 50874 10349 50926
rect 10401 50874 10434 50926
rect 10330 50862 10434 50874
rect 10330 50810 10349 50862
rect 10401 50810 10434 50862
rect 10330 50798 10434 50810
rect 10330 50746 10349 50798
rect 10401 50746 10434 50798
rect 10330 602 10434 50746
<< via2 >>
rect -2933 87645 -1197 87655
rect -2933 87529 -1197 87645
rect -2933 87519 -1197 87529
rect -2005 86130 -1709 86506
rect -1434 85509 -1218 85885
rect 25223 85567 25599 85863
rect 29832 85550 30368 85846
rect -1019 84841 -803 85137
rect 24852 84789 25308 85165
rect 25761 84435 26377 84571
rect -753 81043 -457 81179
rect -2933 77312 -1597 77330
rect -2933 77132 -2931 77312
rect -2931 77132 -1599 77312
rect -1599 77132 -1597 77312
rect -2933 77114 -1597 77132
rect -1024 76938 -328 76948
rect -1024 76822 -1022 76938
rect -1022 76822 -330 76938
rect -330 76822 -328 76938
rect -1024 76812 -328 76822
rect -3100 63574 -2644 63584
rect -3100 63458 -2644 63574
rect -3100 63448 -2644 63458
rect -3105 56371 -2649 56381
rect -3105 56255 -3095 56371
rect -3095 56255 -2659 56371
rect -2659 56255 -2649 56371
rect -3105 56245 -2649 56255
rect -3107 50358 -2651 50368
rect -3107 50242 -3097 50358
rect -3097 50242 -2661 50358
rect -2661 50242 -2651 50358
rect -3107 50232 -2651 50242
rect -3078 43833 -3068 43969
rect -3068 43833 -2632 43969
rect -2632 43833 -2622 43969
rect -3047 36861 -2671 36997
rect -3070 30601 -2614 30619
rect -3070 30421 -2614 30601
rect -3070 30403 -2614 30421
rect -3032 23772 -2656 23782
rect -3032 23656 -3030 23772
rect -3030 23656 -2658 23772
rect -2658 23656 -2656 23772
rect -3032 23646 -2656 23656
rect -3048 16768 -2672 16778
rect -3048 16652 -3046 16768
rect -3046 16652 -2674 16768
rect -2674 16652 -2672 16768
rect -3048 16642 -2672 16652
rect -3030 9978 -2574 9988
rect -3030 9862 -2574 9978
rect -3030 9852 -2574 9862
rect -3004 2773 -2548 2783
rect -3004 2657 -2994 2773
rect -2994 2657 -2558 2773
rect -2558 2657 -2548 2773
rect -3004 2647 -2548 2657
rect 1661 1116 1663 1332
rect 1663 1116 2035 1332
rect 2035 1116 2037 1332
rect 31423 63068 31799 63078
rect 31423 62952 31425 63068
rect 31425 62952 31797 63068
rect 31797 62952 31799 63068
rect 31423 62942 31799 62952
rect 15411 57229 16507 57365
rect 10780 56988 11476 56998
rect 10780 56872 10782 56988
rect 10782 56872 11474 56988
rect 11474 56872 11476 56988
rect 10780 56862 11476 56872
rect 17618 57180 18794 57316
rect 16663 56471 17199 56687
rect 23553 56468 23849 56684
rect 26653 56659 27109 56795
<< metal3 >>
rect 26556 89988 26628 90140
rect 29076 89998 29238 90078
rect 31866 90006 31934 90086
rect 32000 90006 32796 90010
rect 17928 89822 18574 89834
rect 17928 89678 17939 89822
rect 18563 89678 18574 89822
rect 26516 89746 26698 89988
rect 17928 89666 18574 89678
rect 26512 89450 26700 89746
rect 29076 89730 29236 89998
rect 31866 89842 32796 90006
rect 31866 89840 32672 89842
rect 29354 89730 32678 89732
rect 29076 89722 32678 89730
rect 29076 89720 32786 89722
rect 29076 89552 32796 89720
rect 29076 89544 32678 89552
rect 26512 89432 32674 89450
rect 26512 89264 32802 89432
rect 26512 89262 32674 89264
rect -3020 87659 -1118 87692
rect -3020 87515 -2937 87659
rect -1193 87515 -1118 87659
rect -3020 87440 -1118 87515
rect -2096 86511 32490 86542
rect -2096 86506 32046 86511
rect -2096 86130 -2005 86506
rect -1709 86467 32046 86506
rect -1709 86243 17903 86467
rect 18527 86243 32046 86467
rect -1709 86130 32046 86243
rect -2096 86127 32046 86130
rect 32430 86127 32490 86511
rect -2096 86086 32490 86127
rect -2096 85901 32490 85926
rect -2096 85885 31424 85901
rect -2096 85509 -1434 85885
rect -1218 85863 31424 85885
rect -1218 85567 25223 85863
rect 25599 85846 31424 85863
rect 25599 85567 29832 85846
rect -1218 85550 29832 85567
rect 30368 85550 31424 85846
rect -1218 85517 31424 85550
rect 31808 85517 32490 85901
rect -1218 85509 32490 85517
rect -2096 85470 32490 85509
rect -2096 85171 32490 85208
rect -2096 85165 30750 85171
rect -2096 85137 24852 85165
rect -2096 84841 -1019 85137
rect -803 85131 24852 85137
rect -803 84841 21758 85131
rect -2096 84827 21758 84841
rect 21982 84827 24852 85131
rect -2096 84789 24852 84827
rect 25308 84789 30750 85165
rect -2096 84787 30750 84789
rect 31134 84787 32490 85171
rect -2096 84752 32490 84787
rect 25672 84750 26680 84752
rect 25728 84610 26402 84614
rect 25722 84571 32806 84610
rect 25722 84435 25761 84571
rect 26377 84435 32806 84571
rect 25722 84382 32806 84435
rect 25722 84380 32695 84382
rect -3194 81168 -2396 81206
rect -804 81179 -398 81220
rect -804 81168 -753 81179
rect -3194 81050 -753 81168
rect -3194 80996 -2396 81050
rect -804 81043 -753 81050
rect -457 81168 -398 81179
rect -457 81050 -380 81168
rect -457 81043 -398 81050
rect -804 81002 -398 81043
rect -3028 77330 -1522 77362
rect -3028 77294 -2933 77330
rect -1597 77294 -1522 77330
rect -3028 77150 -2937 77294
rect -1593 77150 -1522 77294
rect -3028 77114 -2933 77150
rect -1597 77114 -1522 77150
rect -3028 77088 -1522 77114
rect -3004 77078 -1532 77088
rect -3204 77006 -2404 77008
rect -3204 76994 -1712 77006
rect -3204 76980 -496 76994
rect -3204 76952 -268 76980
rect -3204 76808 -1028 76952
rect -324 76808 -268 76952
rect -3204 76798 -268 76808
rect -2510 76796 -268 76798
rect -2418 76772 -268 76796
rect -1044 76756 -268 76772
rect -10 71091 32464 71154
rect -10 70307 15754 71091
rect 16218 71060 32464 71091
rect 16218 70356 20053 71060
rect 20357 71055 32464 71060
rect 20357 70356 32071 71055
rect 16218 70351 32071 70356
rect 32375 70351 32464 71055
rect 16218 70307 32464 70351
rect -10 70280 32464 70307
rect -10 69912 32085 70010
rect -10 69845 18376 69912
rect -10 69221 267 69845
rect 891 69221 18376 69845
rect -10 69208 18376 69221
rect 19640 69208 32085 69912
rect -10 69136 32085 69208
rect -3138 63608 -2588 63616
rect -3150 63584 -2352 63608
rect -3150 63448 -3100 63584
rect -2644 63448 -2352 63584
rect 31998 63498 32798 63510
rect 26106 63494 32798 63498
rect -3150 63398 -2352 63448
rect 23626 63268 32798 63494
rect 23626 63262 27072 63268
rect 31998 63264 32798 63268
rect 31392 63082 31842 63104
rect 31392 62938 31419 63082
rect 31803 62938 31842 63082
rect 31392 62908 31842 62938
rect 26277 62476 31183 62519
rect 26277 62412 30755 62476
rect 30819 62412 30835 62476
rect 30899 62412 30915 62476
rect 30979 62412 30995 62476
rect 31059 62412 31075 62476
rect 31139 62412 31183 62476
rect 26277 62361 31183 62412
rect 28898 59253 32474 59290
rect 25975 59205 32474 59253
rect 25975 59061 32057 59205
rect 32441 59061 32474 59205
rect 25975 59027 32474 59061
rect 28898 58994 32474 59027
rect 15380 57369 16564 57404
rect 15380 57225 15407 57369
rect 16511 57225 16564 57369
rect 15380 57188 16564 57225
rect 17566 57320 18858 57362
rect 17566 57316 17654 57320
rect 18758 57316 18858 57320
rect 17566 57180 17618 57316
rect 18794 57180 18858 57316
rect 17566 57176 17654 57180
rect 18758 57176 18858 57180
rect 17566 57152 18858 57176
rect 10766 57002 11504 57022
rect 10766 56998 10816 57002
rect 11440 56998 11504 57002
rect 10766 56862 10780 56998
rect 11476 56862 11504 56998
rect 10766 56858 10816 56862
rect 11440 56858 11504 56862
rect 10766 56822 11504 56858
rect 26592 56799 27174 56868
rect 16618 56691 17240 56712
rect 16618 56467 16659 56691
rect 17203 56467 17240 56691
rect 16618 56438 17240 56467
rect 23470 56688 23944 56772
rect 23470 56464 23549 56688
rect 23853 56464 23944 56688
rect 26592 56655 26649 56799
rect 27113 56655 27174 56799
rect 26592 56592 27174 56655
rect -3152 56381 -2354 56416
rect 23470 56400 23944 56464
rect -3152 56245 -3105 56381
rect -2649 56245 -2354 56381
rect -3152 56206 -2354 56245
rect -3208 50368 -2400 50408
rect -3208 50232 -3107 50368
rect -2651 50232 -2400 50368
rect -3208 50194 -2400 50232
rect -3134 50188 -2588 50194
rect -3114 44012 -2584 44020
rect -3206 43969 -2398 44012
rect -3206 43833 -3078 43969
rect -2622 43833 -2398 43969
rect -3206 43798 -2398 43833
rect -3114 43788 -2584 43798
rect -3208 36997 -2398 37054
rect -3208 36861 -3047 36997
rect -2671 36861 -2398 36997
rect -3208 36798 -2398 36861
rect -3122 36794 -2584 36798
rect -3204 30619 -2394 30636
rect -3204 30403 -3070 30619
rect -2614 30403 -2394 30619
rect -3204 30380 -2394 30403
rect -3204 23782 -2394 23844
rect -3204 23646 -3032 23782
rect -2656 23646 -2394 23782
rect -3204 23588 -2394 23646
rect -3210 16778 -2400 16856
rect -3210 16642 -3048 16778
rect -2672 16642 -2400 16778
rect -3210 16600 -2400 16642
rect -3204 9988 -2394 10054
rect -3204 9852 -3030 9988
rect -2574 9852 -2394 9988
rect -3204 9798 -2394 9852
rect 11640 6538 30488 6916
rect 178 6174 382 6428
rect 546 5818 780 6170
rect -3200 3828 -2390 3840
rect -3200 3590 362 3828
rect -3200 3584 -2390 3590
rect -3206 3450 -2396 3462
rect 541 3450 779 3907
rect 11600 3698 30448 4076
rect -3206 3212 779 3450
rect -3206 3206 -2396 3212
rect -3204 2783 -2394 2826
rect -3204 2647 -3004 2783
rect -2548 2647 -2394 2783
rect -3204 2570 -2394 2647
rect 1620 1336 2088 1394
rect 1620 1112 1657 1336
rect 2041 1112 2088 1336
rect 1620 1018 2088 1112
rect 2296 1315 2740 1370
rect 2296 1091 2323 1315
rect 2707 1091 2740 1315
rect 2296 1048 2740 1091
rect 5580 1362 6064 1420
rect 5580 1138 5635 1362
rect 6019 1138 6064 1362
rect 5580 1068 6064 1138
rect 11620 920 30468 1298
rect -3214 392 -2406 394
rect -98 392 32486 396
rect -3214 333 32486 392
rect -3214 109 2329 333
rect 2713 331 32486 333
rect 2713 109 30770 331
rect -3214 107 30770 109
rect 31154 107 32486 331
rect -3214 30 32486 107
rect -3038 24 32486 30
rect -104 20 32486 24
rect -3014 -86 32486 -78
rect -3200 -123 32486 -86
rect -3200 -180 31459 -123
rect -3200 -404 1661 -180
rect 2045 -404 31459 -180
rect -3200 -427 31459 -404
rect 31763 -427 32486 -123
rect -3200 -450 32486 -427
rect -3014 -454 32486 -450
rect -3204 -596 -2396 -594
rect -3204 -643 32486 -596
rect -3204 -700 32073 -643
rect -3204 -924 5629 -700
rect 6013 -924 32073 -700
rect -3204 -947 32073 -924
rect 32377 -947 32486 -643
rect -3204 -958 32486 -947
rect -2992 -972 32486 -958
<< via3 >>
rect 17939 89678 18563 89822
rect -2937 87655 -1193 87659
rect -2937 87519 -2933 87655
rect -2933 87519 -1197 87655
rect -1197 87519 -1193 87655
rect -2937 87515 -1193 87519
rect 17903 86243 18527 86467
rect 32046 86127 32430 86511
rect 31424 85517 31808 85901
rect 21758 84827 21982 85131
rect 30750 84787 31134 85171
rect -2937 77150 -2933 77294
rect -2933 77150 -1597 77294
rect -1597 77150 -1593 77294
rect -1028 76948 -324 76952
rect -1028 76812 -1024 76948
rect -1024 76812 -328 76948
rect -328 76812 -324 76948
rect -1028 76808 -324 76812
rect 15754 70307 16218 71091
rect 20053 70356 20357 71060
rect 32071 70351 32375 71055
rect 267 69221 891 69845
rect 18376 69208 19640 69912
rect 31419 63078 31803 63082
rect 31419 62942 31423 63078
rect 31423 62942 31799 63078
rect 31799 62942 31803 63078
rect 31419 62938 31803 62942
rect 30755 62412 30819 62476
rect 30835 62412 30899 62476
rect 30915 62412 30979 62476
rect 30995 62412 31059 62476
rect 31075 62412 31139 62476
rect 32057 59061 32441 59205
rect 15407 57365 16511 57369
rect 15407 57229 15411 57365
rect 15411 57229 16507 57365
rect 16507 57229 16511 57365
rect 15407 57225 16511 57229
rect 17654 57316 18758 57320
rect 17654 57180 18758 57316
rect 17654 57176 18758 57180
rect 10816 56998 11440 57002
rect 10816 56862 11440 56998
rect 10816 56858 11440 56862
rect 16659 56687 17203 56691
rect 16659 56471 16663 56687
rect 16663 56471 17199 56687
rect 17199 56471 17203 56687
rect 16659 56467 17203 56471
rect 23549 56684 23853 56688
rect 23549 56468 23553 56684
rect 23553 56468 23849 56684
rect 23849 56468 23853 56684
rect 23549 56464 23853 56468
rect 26649 56795 27113 56799
rect 26649 56659 26653 56795
rect 26653 56659 27109 56795
rect 27109 56659 27113 56795
rect 26649 56655 27113 56659
rect 1657 1332 2041 1336
rect 1657 1116 1661 1332
rect 1661 1116 2037 1332
rect 2037 1116 2041 1332
rect 1657 1112 2041 1116
rect 2323 1091 2707 1315
rect 5635 1138 6019 1362
rect 2329 109 2713 333
rect 30770 107 31154 331
rect 1661 -404 2045 -180
rect 31459 -427 31763 -123
rect 5629 -924 6013 -700
rect 32073 -947 32377 -643
<< metal4 >>
rect 17888 89864 18638 89874
rect 17826 89822 18638 89864
rect 17826 89678 17939 89822
rect 18563 89678 18638 89822
rect 17826 89630 18638 89678
rect -2972 87692 -2664 87694
rect -3020 87659 -1118 87692
rect -3020 87515 -2937 87659
rect -1193 87515 -1118 87659
rect -3020 87440 -1118 87515
rect -2972 77362 -2664 87440
rect 17826 86467 18616 89630
rect 17826 86243 17903 86467
rect 18527 86243 18616 86467
rect 17826 86122 18616 86243
rect 21710 85131 22052 90966
rect 21710 84827 21758 85131
rect 21982 84827 22052 85131
rect 21710 84742 22052 84827
rect 30726 85171 31182 86542
rect 30726 84787 30750 85171
rect 31134 84787 31182 85171
rect -3028 77294 -1522 77362
rect -3028 77150 -2937 77294
rect -1593 77150 -1522 77294
rect -3028 77088 -1522 77150
rect -3004 77078 -1532 77088
rect -1020 76982 -888 76984
rect -1020 76980 -802 76982
rect -1044 76952 -268 76980
rect -1044 76808 -1028 76952
rect -324 76808 -268 76952
rect -1044 76756 -268 76808
rect -1020 57056 -802 76756
rect 205 69845 954 82386
rect 19528 76550 19938 76558
rect 19292 76536 19938 76550
rect 19292 75334 20456 76536
rect 19292 75170 19938 75334
rect 205 69221 267 69845
rect 891 69221 954 69845
rect 205 69136 954 69221
rect 15708 71091 16282 71166
rect 15708 70307 15754 71091
rect 16218 70307 16282 71091
rect 15708 57404 16282 70307
rect 19295 70034 19705 75170
rect 19980 74248 20444 74268
rect 19980 73046 20466 74248
rect 19980 72664 20444 73046
rect 19980 71060 20438 72664
rect 19980 70356 20053 71060
rect 20357 70356 20438 71060
rect 19980 70306 20438 70356
rect 18300 69912 19705 70034
rect 18300 69208 18376 69912
rect 19640 69208 19705 69912
rect 18300 69143 19705 69208
rect 18300 69140 19682 69143
rect 15380 57369 16564 57404
rect 15380 57225 15407 57369
rect 16511 57225 16564 57369
rect 18314 57362 18986 69140
rect 15380 57188 16564 57225
rect 17566 57320 18986 57362
rect -1018 57032 -802 57056
rect 17566 57176 17654 57320
rect 18758 57176 18986 57320
rect 17566 57164 18986 57176
rect 30726 62476 31182 84787
rect 30726 62412 30755 62476
rect 30819 62412 30835 62476
rect 30899 62412 30915 62476
rect 30979 62412 30995 62476
rect 31059 62412 31075 62476
rect 31139 62412 31182 62476
rect 17566 57152 18858 57164
rect -1018 57022 11482 57032
rect -1018 57002 11504 57022
rect -1018 56858 10816 57002
rect 11440 56858 11504 57002
rect -1018 56822 11504 56858
rect -1018 56816 11482 56822
rect 16614 56712 17238 56740
rect 16614 56699 17240 56712
rect 16614 56463 16652 56699
rect 16888 56691 16972 56699
rect 16888 56463 16972 56467
rect 17208 56463 17240 56699
rect 16614 56440 17240 56463
rect 16618 56438 17240 56440
rect 17566 56222 18376 57152
rect 26592 56865 27174 56868
rect 26592 56799 26763 56865
rect 26999 56799 27174 56865
rect 23470 56697 23944 56772
rect 23470 56688 23584 56697
rect 23820 56688 23944 56697
rect 23470 56464 23549 56688
rect 23853 56464 23944 56688
rect 26592 56655 26649 56799
rect 27113 56655 27174 56799
rect 26592 56629 26763 56655
rect 26999 56629 27174 56655
rect 26592 56592 27174 56629
rect 23470 56461 23584 56464
rect 23820 56461 23944 56464
rect 23470 56400 23944 56461
rect 1624 1336 2092 1370
rect 5584 1362 6064 1420
rect 1624 1112 1657 1336
rect 2041 1112 2092 1336
rect 1624 -180 2092 1112
rect 2292 1315 2744 1354
rect 2292 1091 2323 1315
rect 2707 1091 2744 1315
rect 2292 333 2744 1091
rect 2292 109 2329 333
rect 2713 109 2744 333
rect 2292 30 2744 109
rect 5584 1138 5635 1362
rect 6019 1138 6064 1362
rect 1624 -404 1661 -180
rect 2045 -404 2092 -180
rect 1624 -454 2092 -404
rect 5584 -700 6064 1138
rect 12493 768 12927 9651
rect 14894 768 15338 9634
rect 17188 768 17632 9622
rect 19618 768 20062 9602
rect 21976 768 22420 9654
rect 24364 768 24808 9622
rect 26834 768 27278 9588
rect 29192 768 29636 9622
rect 5584 -924 5629 -700
rect 6013 -924 6064 -700
rect 5584 -982 6064 -924
rect 30726 331 31182 62412
rect 31388 85901 31844 86548
rect 31388 85517 31424 85901
rect 31808 85517 31844 85901
rect 31388 63082 31844 85517
rect 31388 62938 31419 63082
rect 31803 62938 31844 63082
rect 31388 1412 31844 62938
rect 30726 107 30770 331
rect 31154 107 31182 331
rect 30726 -992 31182 107
rect 31382 32 31844 1412
rect 31388 -123 31844 32
rect 31388 -427 31459 -123
rect 31763 -427 31844 -123
rect 31388 -992 31844 -427
rect 32018 86511 32474 86536
rect 32018 86127 32046 86511
rect 32430 86127 32474 86511
rect 32018 71055 32474 86127
rect 32018 70351 32071 71055
rect 32375 70351 32474 71055
rect 32018 59205 32474 70351
rect 32018 59061 32057 59205
rect 32441 59061 32474 59205
rect 32018 1102 32474 59061
rect 32018 -278 32480 1102
rect 32018 -643 32474 -278
rect 32018 -947 32073 -643
rect 32377 -947 32474 -643
rect 32018 -992 32474 -947
<< via4 >>
rect 16652 56691 16888 56699
rect 16972 56691 17208 56699
rect 16652 56467 16659 56691
rect 16659 56467 16888 56691
rect 16972 56467 17203 56691
rect 17203 56467 17208 56691
rect 16652 56463 16888 56467
rect 16972 56463 17208 56467
rect 26763 56799 26999 56865
rect 23584 56688 23820 56697
rect 23584 56464 23820 56688
rect 26763 56655 26999 56799
rect 26763 56629 26999 56655
rect 23584 56461 23820 56464
<< metal5 >>
rect 26588 56914 27172 56916
rect 26586 56865 27174 56914
rect 16612 56752 17244 56764
rect 23470 56752 23944 56772
rect 16450 56699 23944 56752
rect 16450 56463 16652 56699
rect 16888 56463 16972 56699
rect 17208 56697 23944 56699
rect 17208 56463 23584 56697
rect 16450 56461 23584 56463
rect 23820 56461 23944 56697
rect 26586 56629 26763 56865
rect 26999 56629 27174 56865
rect 26586 56592 27174 56629
rect 26588 56590 27172 56592
rect 16450 56416 23944 56461
rect 16618 39048 17242 56416
rect 23470 56400 23944 56416
rect 16618 38424 19976 39048
rect 26710 30424 27170 56590
rect 19502 29964 27170 30424
use EF_AMUX21_ARRAY  EF_AMUX21_ARRAY_0
timestamp 1694077897
transform 0 1 978 -1 0 20186
box -48698 -806 19118 7110
use EF_AMUX0801  EF_AMUX0801_0
timestamp 1694077897
transform 1 0 -5031 0 -1 94698
box 3148 -1716 37700 7264
use EF_BANK_CAP_10  EF_BANK_CAP_10_0
timestamp 1694077897
transform 1 0 18760 0 1 43012
box -7958 -33880 11700 13322
use EF_BUF3V3  EF_BUF3V3_0
timestamp 1694077897
transform 0 -1 17605 1 0 61545
box -4547 -3901 2817 6641
use EF_R2RVC  EF_R2RVC_0
timestamp 1694077897
transform 0 -1 30236 1 0 72561
box -200 -265 11765 10234
use EF_SW_RST  EF_SW_RST_1
timestamp 1694077897
transform 1 0 27330 0 -1 63109
box -4247 -398 2232 6031
use sample_and_hold  sample_and_hold_0
timestamp 1694077897
transform 1 0 -652 0 1 72114
box 0 -114 19469 11183
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_0
timestamp 1694077897
transform 0 1 29442 -1 0 7716
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_1
timestamp 1694077897
transform 0 1 29438 -1 0 2096
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_2
timestamp 1694077897
transform 0 1 15040 -1 0 7676
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_3
timestamp 1694077897
transform 0 1 17444 -1 0 7688
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_4
timestamp 1694077897
transform 0 1 19844 -1 0 7702
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_5
timestamp 1694077897
transform 0 1 12638 -1 0 7672
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_6
timestamp 1694077897
transform 0 1 29462 -1 0 4906
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_7
timestamp 1694077897
transform 0 1 22246 -1 0 7702
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_8
timestamp 1694077897
transform 0 1 24650 -1 0 7702
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_9
timestamp 1694077897
transform 0 1 27056 -1 0 7702
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_10
timestamp 1694077897
transform 0 1 12644 -1 0 4880
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_11
timestamp 1694077897
transform 0 1 15058 -1 0 4892
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_12
timestamp 1694077897
transform 0 1 17456 -1 0 4892
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_13
timestamp 1694077897
transform 0 1 19862 -1 0 4896
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_14
timestamp 1694077897
transform 0 1 22260 -1 0 4902
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_15
timestamp 1694077897
transform 0 1 24662 -1 0 4916
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_16
timestamp 1694077897
transform 0 1 27060 -1 0 4912
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_17
timestamp 1694077897
transform 0 1 12642 -1 0 2086
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_18
timestamp 1694077897
transform 0 1 15044 -1 0 2086
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_19
timestamp 1694077897
transform 0 1 17446 -1 0 2106
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_20
timestamp 1694077897
transform 0 1 19852 -1 0 2086
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_21
timestamp 1694077897
transform 0 1 22240 -1 0 2096
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_22
timestamp 1694077897
transform 0 1 24638 -1 0 2086
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB#0  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_23
timestamp 1694077897
transform 0 1 27040 -1 0 2100
box -1186 -1040 1186 1040
<< labels >>
flabel metal2 s 27104 72785 27104 72785 0 FreeSans 661 270 0 0 VINM
flabel metal3 s 19214 69388 19496 69666 0 FreeSans 1025 0 0 0 VSS
port 1 nsew
flabel metal3 s -3194 80996 -2396 81206 0 FreeSans 2500 0 0 0 HOLD
port 2 nsew
flabel metal3 s -3202 76798 -2404 77008 0 FreeSans 2500 0 0 0 EN
port 3 nsew
flabel metal3 s -3150 63398 -2352 63608 0 FreeSans 2500 0 0 0 DATA[9]
port 4 nsew
flabel metal3 s -3152 56206 -2354 56416 0 FreeSans 2500 0 0 0 DATA[8]
port 5 nsew
flabel metal3 s -3208 50194 -2400 50408 0 FreeSans 2500 0 0 0 DATA[7]
port 6 nsew
flabel metal3 s -3206 43798 -2398 44012 0 FreeSans 2500 0 0 0 DATA[6]
port 7 nsew
flabel metal3 s -3208 36798 -2398 37054 0 FreeSans 2500 0 0 0 DATA[5]
port 8 nsew
flabel metal3 s -3204 30380 -2394 30636 0 FreeSans 2500 0 0 0 DATA[4]
port 9 nsew
flabel metal3 s -3204 23588 -2394 23844 0 FreeSans 2500 0 0 0 DATA[3]
port 10 nsew
flabel metal3 s -3210 16600 -2400 16856 0 FreeSans 2500 0 0 0 DATA[2]
port 11 nsew
flabel metal3 s -3204 9798 -2394 10054 0 FreeSans 2500 0 0 0 DATA[1]
port 12 nsew
flabel metal3 s -3200 3584 -2390 3840 0 FreeSans 2500 0 0 0 VL
port 13 nsew
flabel metal3 s -3206 3206 -2396 3462 0 FreeSans 2500 0 0 0 VH
port 14 nsew
flabel metal3 s -3204 2570 -2394 2826 0 FreeSans 2500 0 0 0 DATA[0]
port 15 nsew
flabel metal3 s -3214 30 -2406 394 0 FreeSans 2500 0 0 0 DVDD
port 16 nsew
flabel metal3 s -3200 -450 -2392 -86 0 FreeSans 2500 0 0 0 DVSS
port 17 nsew
flabel metal3 s -3204 -958 -2396 -594 0 FreeSans 2500 0 0 0 VDD
port 18 nsew
flabel metal3 s 32000 89842 32796 90010 0 FreeSans 2500 0 0 0 B[0]
port 19 nsew
flabel metal3 s 32000 89552 32796 89720 0 FreeSans 2500 0 0 0 B[1]
port 20 nsew
flabel metal3 s 32006 89264 32802 89432 0 FreeSans 2500 0 0 0 B[2]
port 21 nsew
flabel metal3 s 31956 84382 32806 84610 0 FreeSans 2500 0 0 0 CMP
port 22 nsew
flabel metal3 s 31998 63264 32798 63510 0 FreeSans 2500 0 0 0 RST
port 23 nsew
flabel metal2 s 1152 95998 1346 96802 0 FreeSans 2000 0 0 0 VIN[7]
port 24 nsew
flabel metal2 s 4582 95818 4794 96806 0 FreeSans 2000 0 0 0 VIN[6]
port 25 nsew
flabel metal2 s 7924 95818 8136 96806 0 FreeSans 2000 0 0 0 VIN[5]
port 26 nsew
flabel metal2 s 11350 95812 11562 96800 0 FreeSans 2000 0 0 0 VIN[4]
port 27 nsew
flabel metal2 s 14700 95818 14912 96806 0 FreeSans 2000 0 0 0 VIN[3]
port 28 nsew
flabel metal2 s 18178 95826 18390 96814 0 FreeSans 2000 0 0 0 VIN[2]
port 29 nsew
flabel metal2 s 21494 95818 21706 96806 0 FreeSans 2000 0 0 0 VIN[1]
port 30 nsew
flabel metal2 s 24870 95818 25082 96806 0 FreeSans 2000 0 0 0 VIN[0]
port 31 nsew
<< end >>
