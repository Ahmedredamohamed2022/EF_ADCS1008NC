magic
tech sky130A
magscale 1 2
timestamp 1699926577
<< metal1 >>
rect 174 5490 312 5888
rect 2612 2920 2804 3244
rect 2876 776 3068 2312
rect 252 705 590 718
rect 252 589 271 705
rect 579 589 590 705
rect 252 576 590 589
rect 1854 710 2164 716
rect 1854 594 1887 710
rect 2131 594 2164 710
rect 2816 698 3070 776
rect 2876 692 3068 698
rect 1854 582 2164 594
rect 348 326 598 530
<< via1 >>
rect 271 589 579 705
rect 1887 594 2131 710
<< metal2 >>
rect 158 4083 822 4102
rect 158 3947 182 4083
rect 798 3947 822 4083
rect 158 3928 822 3947
rect 56 1338 228 2354
rect 790 1159 1296 1188
rect 790 1103 815 1159
rect 871 1103 895 1159
rect 951 1103 975 1159
rect 1031 1103 1055 1159
rect 1111 1103 1135 1159
rect 1191 1103 1215 1159
rect 1271 1103 1296 1159
rect 790 1074 1296 1103
rect 260 705 590 718
rect 260 589 271 705
rect 579 589 590 705
rect 260 576 590 589
rect 1854 710 2164 716
rect 1854 594 1887 710
rect 2131 594 2164 710
rect 1854 582 2164 594
<< via2 >>
rect 182 3947 798 4083
rect 815 1103 871 1159
rect 895 1103 951 1159
rect 975 1103 1031 1159
rect 1055 1103 1111 1159
rect 1135 1103 1191 1159
rect 1215 1103 1271 1159
rect 277 619 333 675
rect 357 619 413 675
rect 437 619 493 675
rect 517 619 573 675
rect 1905 627 1961 683
rect 1985 627 2041 683
rect 2065 627 2121 683
<< metal3 >>
rect 80 4083 1940 4128
rect 80 3947 182 4083
rect 798 3947 1940 4083
rect 80 3904 1940 3947
rect 90 3902 1940 3904
rect 758 1159 1358 3902
rect 758 1103 815 1159
rect 871 1103 895 1159
rect 951 1103 975 1159
rect 1031 1103 1055 1159
rect 1111 1103 1135 1159
rect 1191 1103 1215 1159
rect 1271 1103 1358 1159
rect 758 1026 1358 1103
rect 52 683 2188 736
rect 52 675 1905 683
rect 52 619 277 675
rect 333 619 357 675
rect 413 619 437 675
rect 493 619 517 675
rect 573 627 1905 675
rect 1961 627 1985 683
rect 2041 627 2065 683
rect 2121 627 2188 683
rect 573 619 2188 627
rect 52 578 2188 619
rect 260 576 590 578
use array_1lsm  array_1lsm_0
timestamp 1699926577
transform 1 0 -2700 0 1 -202
box 2700 202 5594 1958
use array_1tgm  array_1tgm_0
timestamp 1699926577
transform -1 0 4964 0 1 1916
box 1896 0 4886 4141
<< labels >>
flabel metal1 s 2700 3074 2742 3132 0 FreeSans 625 0 0 0 in0
port 1 nsew
flabel metal1 s 436 344 454 354 0 FreeSans 625 0 0 0 l0
port 2 nsew
flabel metal2 s 108 1952 124 1970 0 FreeSans 506 0 0 0 vss
port 3 nsew
flabel metal1 s 238 5644 260 5726 0 FreeSans 506 0 0 0 vo
port 4 nsew
flabel metal3 s 104 3976 124 4042 0 FreeSans 506 0 0 0 vdd3p3
port 5 nsew
flabel metal3 s 1020 598 1032 616 0 FreeSans 506 0 0 0 vdd1p8
port 6 nsew
<< end >>
