magic
tech sky130A
magscale 1 2
timestamp 1699926577
<< metal1 >>
rect -3990 5720 -3796 5998
rect -690 5738 -494 6004
rect -1512 3180 -1374 3198
rect -1512 1976 -1501 3180
rect -1385 1976 -1374 3180
rect -1512 1958 -1374 1976
rect 1782 3196 1942 3202
rect 1782 1928 1804 3196
rect 1920 1928 1942 3196
rect 1782 1922 1942 1928
rect -3836 498 -3560 548
rect -3836 382 -3815 498
rect -3571 382 -3560 498
rect -3836 332 -3560 382
rect -524 499 -242 544
rect -524 383 -477 499
rect -297 383 -242 499
rect -524 334 -242 383
rect -1458 196 1300 208
rect -1496 170 1300 196
rect -1496 54 -1485 170
rect -1241 54 1300 170
rect -1496 28 1300 54
rect 1798 163 1934 172
rect 1798 47 1808 163
rect 1924 47 1934 163
rect 1798 38 1934 47
rect -1458 12 1300 28
<< via1 >>
rect -1501 1976 -1385 3180
rect 1804 1928 1920 3196
rect -3815 382 -3571 498
rect -477 383 -297 499
rect -1485 54 -1241 170
rect 1808 47 1924 163
<< metal2 >>
rect -1532 3180 -1348 3228
rect -1532 3166 -1501 3180
rect -1385 3166 -1348 3180
rect -1532 1990 -1511 3166
rect -1375 1990 -1348 3166
rect -1532 1976 -1501 1990
rect -1385 1976 -1348 1990
rect -1532 1908 -1348 1976
rect 1766 3196 1956 3224
rect 1766 3190 1804 3196
rect 1920 3190 1956 3196
rect 1766 1934 1794 3190
rect 1930 1934 1956 3190
rect 1766 1928 1804 1934
rect 1920 1928 1956 1934
rect 1766 1896 1956 1928
rect -3836 498 -3560 548
rect -524 542 -242 544
rect -3836 382 -3815 498
rect -3571 382 -3560 498
rect -3836 332 -3560 382
rect -526 499 -242 542
rect -526 383 -477 499
rect -297 383 -242 499
rect -526 334 -242 383
rect -3790 -150 -3576 332
rect -1524 180 -1206 206
rect -1524 170 -1471 180
rect -1255 170 -1206 180
rect -1524 54 -1485 170
rect -1241 54 -1206 170
rect -1524 44 -1471 54
rect -1255 44 -1206 54
rect -1524 8 -1206 44
rect -3792 -210 -3238 -150
rect -3792 -346 -3743 -210
rect -3287 -346 -3238 -210
rect -3792 -396 -3238 -346
rect -526 -194 -246 334
rect 1774 163 1954 192
rect 1774 133 1808 163
rect 1924 133 1954 163
rect 1774 77 1798 133
rect 1934 77 1954 133
rect 1774 47 1808 77
rect 1924 47 1954 77
rect 1774 12 1954 47
rect -526 -228 -242 -194
rect -526 -364 -486 -228
rect -270 -364 -242 -228
rect -526 -398 -242 -364
<< via2 >>
rect -1511 1990 -1501 3166
rect -1501 1990 -1385 3166
rect -1385 1990 -1375 3166
rect 1794 1934 1804 3190
rect 1804 1934 1920 3190
rect 1920 1934 1930 3190
rect -1471 170 -1255 180
rect -1471 54 -1255 170
rect -1471 44 -1255 54
rect -3743 -346 -3287 -210
rect 1798 77 1808 133
rect 1808 77 1854 133
rect 1878 77 1924 133
rect 1924 77 1934 133
rect -486 -364 -270 -228
<< metal3 >>
rect -2505 3856 191 4082
rect -1532 3170 -1348 3228
rect -1532 3166 -1475 3170
rect -1411 3166 -1348 3170
rect -1532 1990 -1511 3166
rect -1375 1990 -1348 3166
rect -1532 1986 -1475 1990
rect -1411 1986 -1348 1990
rect -1532 1908 -1348 1986
rect 1766 3194 1956 3224
rect 1766 1930 1790 3194
rect 1934 1930 1956 3194
rect 1766 1896 1956 1930
rect -2081 590 345 748
rect -1524 184 -1206 206
rect -1524 40 -1475 184
rect -1251 40 -1206 184
rect -1524 8 -1206 40
rect 1774 137 1954 192
rect 1774 133 1834 137
rect 1898 133 1954 137
rect 1774 77 1798 133
rect 1934 77 1954 133
rect 1774 73 1834 77
rect 1898 73 1954 77
rect 1774 12 1954 73
rect -3660 -150 -3238 -148
rect -3792 -194 -3238 -150
rect -3792 -210 -242 -194
rect -3792 -346 -3743 -210
rect -3287 -228 -242 -210
rect -3287 -346 -486 -228
rect -3792 -364 -486 -346
rect -270 -364 -242 -228
rect -3792 -394 -242 -364
rect -3792 -396 -3238 -394
<< via3 >>
rect -1475 3166 -1411 3170
rect -1475 3106 -1411 3166
rect -1475 3026 -1411 3090
rect -1475 2946 -1411 3010
rect -1475 2866 -1411 2930
rect -1475 2786 -1411 2850
rect -1475 2706 -1411 2770
rect -1475 2626 -1411 2690
rect -1475 2546 -1411 2610
rect -1475 2466 -1411 2530
rect -1475 2386 -1411 2450
rect -1475 2306 -1411 2370
rect -1475 2226 -1411 2290
rect -1475 2146 -1411 2210
rect -1475 2066 -1411 2130
rect -1475 1990 -1411 2050
rect -1475 1986 -1411 1990
rect 1790 3190 1934 3194
rect 1790 1934 1794 3190
rect 1794 1934 1930 3190
rect 1930 1934 1934 3190
rect 1790 1930 1934 1934
rect -1475 180 -1251 184
rect -1475 44 -1471 180
rect -1471 44 -1255 180
rect -1255 44 -1251 180
rect -1475 40 -1251 44
rect 1834 133 1898 137
rect 1834 77 1854 133
rect 1854 77 1878 133
rect 1878 77 1898 133
rect 1834 73 1898 77
<< metal4 >>
rect -1532 3170 -1348 3228
rect -1532 3106 -1475 3170
rect -1411 3106 -1348 3170
rect -1532 3090 -1348 3106
rect -1532 3026 -1475 3090
rect -1411 3026 -1348 3090
rect -1532 3010 -1348 3026
rect -1532 2946 -1475 3010
rect -1411 2946 -1348 3010
rect -1532 2930 -1348 2946
rect -1532 2866 -1475 2930
rect -1411 2866 -1348 2930
rect -1532 2850 -1348 2866
rect -1532 2786 -1475 2850
rect -1411 2786 -1348 2850
rect -1532 2770 -1348 2786
rect -1532 2706 -1475 2770
rect -1411 2706 -1348 2770
rect -1532 2690 -1348 2706
rect -1532 2626 -1475 2690
rect -1411 2626 -1348 2690
rect -1532 2610 -1348 2626
rect -1532 2546 -1475 2610
rect -1411 2546 -1348 2610
rect -1532 2530 -1348 2546
rect -1532 2466 -1475 2530
rect -1411 2466 -1348 2530
rect -1532 2450 -1348 2466
rect -1532 2386 -1475 2450
rect -1411 2386 -1348 2450
rect -1532 2370 -1348 2386
rect -1532 2306 -1475 2370
rect -1411 2306 -1348 2370
rect -1532 2290 -1348 2306
rect -1532 2226 -1475 2290
rect -1411 2226 -1348 2290
rect -1532 2210 -1348 2226
rect -1532 2146 -1475 2210
rect -1411 2146 -1348 2210
rect -1532 2130 -1348 2146
rect -1532 2066 -1475 2130
rect -1411 2066 -1348 2130
rect -1532 2050 -1348 2066
rect -1532 1986 -1475 2050
rect -1411 1986 -1348 2050
rect -1532 1908 -1348 1986
rect -1524 206 -1348 1908
rect 1766 3194 1956 3224
rect 1766 1930 1790 3194
rect 1934 1930 1956 3194
rect 1766 1896 1956 1930
rect -1524 184 -1206 206
rect -1524 40 -1475 184
rect -1251 40 -1206 184
rect -1524 8 -1206 40
rect 1774 137 1954 1896
rect 1774 73 1834 137
rect 1898 73 1954 137
rect 1774 12 1954 73
use array_1ls_1tgm  array_1ls_1tgm_0
timestamp 1699926577
transform 1 0 -854 0 1 12
box -1539 -257 3674 6057
use array_1ls_1tgm  array_1ls_1tgm_1
timestamp 1699926577
transform 1 0 -4150 0 1 14
box -1539 -257 3674 6057
<< labels >>
flabel metal3 s -1352 3964 -1282 4044 0 FreeSans 3283 0 0 0 VDD
port 1 nsew
flabel metal3 s -1042 616 -974 682 0 FreeSans 3283 0 0 0 DVDD
port 2 nsew
flabel metal1 s -1048 68 -982 122 0 FreeSans 3283 0 0 0 VSS
port 3 nsew
flabel metal3 s -2128 -314 -1996 -226 0 FreeSans 3283 0 0 0 RST
port 4 nsew
flabel metal1 s -628 5816 -596 5880 0 FreeSans 3283 0 0 0 VP1
port 5 nsew
flabel metal1 s -3930 5810 -3880 5882 0 FreeSans 5250 0 0 0 VP2
port 6 nsew
<< end >>
