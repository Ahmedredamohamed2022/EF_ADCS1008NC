magic
tech sky130A
magscale 1 2
timestamp 1699926577
<< locali >>
rect 392 8914 616 9238
rect 940 9202 2054 9238
rect 940 8952 1174 9202
rect 2000 8952 2054 9202
rect 940 8914 2054 8952
rect 392 8734 426 8914
rect 2020 8732 2054 8914
rect 722 8603 830 8646
rect 722 8569 762 8603
rect 796 8569 830 8603
rect 722 8531 830 8569
rect 722 8497 762 8531
rect 796 8497 830 8531
rect 722 8459 830 8497
rect 722 8425 762 8459
rect 796 8425 830 8459
rect 722 8387 830 8425
rect 722 8353 762 8387
rect 796 8353 830 8387
rect 722 8315 830 8353
rect 722 8281 762 8315
rect 796 8281 830 8315
rect 722 8214 830 8281
rect 1692 6610 1778 6648
rect 1428 6585 1778 6610
rect 1428 6551 1441 6585
rect 1475 6551 1513 6585
rect 1547 6551 1585 6585
rect 1619 6551 1657 6585
rect 1691 6551 1729 6585
rect 1763 6551 1778 6585
rect 1428 6524 1778 6551
<< viali >>
rect 1174 8952 2000 9202
rect 762 8569 796 8603
rect 762 8497 796 8531
rect 762 8425 796 8459
rect 762 8353 796 8387
rect 762 8281 796 8315
rect 1441 6551 1475 6585
rect 1513 6551 1547 6585
rect 1585 6551 1619 6585
rect 1657 6551 1691 6585
rect 1729 6551 1763 6585
<< metal1 >>
rect 11011 11152 11403 11182
rect 11011 10908 11052 11152
rect 11360 10908 11403 11152
rect 11011 10151 11403 10908
rect 0 9612 1070 9952
rect 0 9040 200 9101
rect 0 8950 815 9040
rect 0 8901 200 8950
rect 743 8632 815 8950
rect 1013 8655 1070 9612
rect 11011 9267 11021 10151
rect 11393 9267 11403 10151
rect 1118 9202 2060 9238
rect 1118 8952 1174 9202
rect 2000 8952 2060 9202
rect 1118 8914 2060 8952
rect 1912 8702 1986 8914
rect 2014 8738 2060 8914
rect 2014 8702 2020 8738
rect 2054 8702 2060 8738
rect 732 8603 826 8632
rect 732 8569 762 8603
rect 796 8569 826 8603
rect 732 8531 826 8569
rect 732 8497 762 8531
rect 796 8497 826 8531
rect 732 8459 826 8497
rect 732 8425 762 8459
rect 796 8425 826 8459
rect 732 8387 826 8425
rect 732 8353 762 8387
rect 796 8353 826 8387
rect 732 8315 826 8353
rect 732 8281 762 8315
rect 796 8281 826 8315
rect 732 8246 826 8281
rect 386 6474 432 6652
rect 460 6474 534 6652
rect 0 6436 1040 6474
rect 0 6192 830 6436
rect 1010 6192 1040 6436
rect 0 6152 1040 6192
rect 1098 6082 1172 6700
rect 1200 6082 1246 6646
rect 1274 6082 1348 6700
rect 1428 6594 1778 6610
rect 1428 6585 1448 6594
rect 1428 6551 1441 6585
rect 1428 6542 1448 6551
rect 1500 6542 1512 6594
rect 1564 6542 1576 6594
rect 1628 6542 1640 6594
rect 1692 6542 1704 6594
rect 1756 6585 1778 6594
rect 1763 6551 1778 6585
rect 1756 6542 1778 6551
rect 1428 6524 1778 6542
rect 1912 6476 1986 6640
rect 2014 6476 2060 6640
rect 1406 6438 2060 6476
rect 1406 6194 1429 6438
rect 1609 6194 2060 6438
rect 1406 6152 2060 6194
rect 11011 6302 11403 9267
rect 1098 6015 1348 6082
rect 0 5995 3424 6015
rect 0 5303 2543 5995
rect 3363 5303 3424 5995
rect 11011 5994 11054 6302
rect 11362 5994 11403 6302
rect 11011 5949 11403 5994
rect 10725 5488 12368 5842
rect 0 5284 3424 5303
rect 11011 5315 11403 5360
rect 0 4986 3717 5186
rect 11011 5007 11053 5315
rect 11361 5007 11403 5315
rect 0 4831 3717 4841
rect 0 4651 1916 4831
rect 2352 4651 3717 4831
rect 0 4641 3717 4651
rect 11011 4436 11403 5007
rect 11011 4064 11021 4436
rect 11393 4064 11403 4436
rect 2404 2703 3517 2719
rect 2404 2459 2543 2703
rect 3363 2459 3517 2703
rect 2404 2443 3517 2459
rect 2924 1925 3657 2298
rect 11011 2268 11403 4064
rect 2416 1647 2693 1847
rect 2493 1573 2693 1647
rect 2493 1457 2503 1573
rect 2683 1457 2693 1573
rect 2493 1427 2693 1457
rect 2924 1256 3506 1925
rect 2924 941 2963 1256
rect 872 913 1589 929
rect 872 733 884 913
rect 1576 733 1589 913
rect 872 718 1589 733
rect 2402 756 2963 941
rect 3463 756 3506 1256
rect 2402 706 3506 756
rect 11011 680 11021 2268
rect 11393 680 11403 2268
rect 11011 627 11403 680
rect 11546 4996 12150 5196
rect 11546 281 11746 4996
rect 11875 4651 12150 4851
rect 11875 483 11987 4651
rect 19130 4570 19469 4770
rect 11875 452 12216 483
rect 11875 400 11891 452
rect 11943 400 11955 452
rect 12007 400 12019 452
rect 12071 400 12083 452
rect 12135 400 12147 452
rect 12199 400 12216 452
rect 11875 370 12216 400
rect 2478 238 3021 281
rect 2478 -70 2534 238
rect 2970 -70 3021 238
rect 2478 -114 3021 -70
rect 11278 238 11821 281
rect 11278 -70 11334 238
rect 11770 -70 11821 238
rect 11278 -114 11821 -70
<< via1 >>
rect 11052 10908 11360 11152
rect 11021 9267 11393 10151
rect 830 6192 1010 6436
rect 1448 6585 1500 6594
rect 1448 6551 1475 6585
rect 1475 6551 1500 6585
rect 1448 6542 1500 6551
rect 1512 6585 1564 6594
rect 1512 6551 1513 6585
rect 1513 6551 1547 6585
rect 1547 6551 1564 6585
rect 1512 6542 1564 6551
rect 1576 6585 1628 6594
rect 1576 6551 1585 6585
rect 1585 6551 1619 6585
rect 1619 6551 1628 6585
rect 1576 6542 1628 6551
rect 1640 6585 1692 6594
rect 1640 6551 1657 6585
rect 1657 6551 1691 6585
rect 1691 6551 1692 6585
rect 1640 6542 1692 6551
rect 1704 6585 1756 6594
rect 1704 6551 1729 6585
rect 1729 6551 1756 6585
rect 1704 6542 1756 6551
rect 1429 6194 1609 6438
rect 2543 5303 3363 5995
rect 11054 5994 11362 6302
rect 11053 5007 11361 5315
rect 1916 4651 2352 4831
rect 11021 4064 11393 4436
rect 2543 2459 3363 2703
rect 2503 1457 2683 1573
rect 884 733 1576 913
rect 2963 756 3463 1256
rect 11021 680 11393 2268
rect 11891 400 11943 452
rect 11955 400 12007 452
rect 12019 400 12071 452
rect 12083 400 12135 452
rect 12147 400 12199 452
rect 2534 -70 2970 238
rect 11334 -70 11770 238
<< metal2 >>
rect 11011 11152 11403 11182
rect 2515 10932 3391 11027
rect 2515 10710 3685 10932
rect 10732 10756 10958 10932
rect 11011 10908 11052 11152
rect 11360 10908 11403 11152
rect 11011 10836 11403 10908
rect 11477 10756 12149 10942
rect 10732 10710 12149 10756
rect 1428 6594 1778 6610
rect 1428 6542 1448 6594
rect 1500 6542 1512 6594
rect 1564 6542 1576 6594
rect 1628 6542 1640 6594
rect 1692 6542 1704 6594
rect 1756 6542 1778 6594
rect 1428 6524 1778 6542
rect 798 6438 1630 6474
rect 798 6436 1429 6438
rect 798 6192 830 6436
rect 1010 6194 1429 6436
rect 1609 6194 1630 6438
rect 1010 6192 1630 6194
rect 798 6152 1630 6192
rect 1692 3414 1778 6524
rect 2515 5995 3391 10710
rect 10835 10479 11721 10710
rect 2515 5303 2543 5995
rect 3363 5842 3391 5995
rect 11011 10151 11403 10231
rect 11011 9267 11021 10151
rect 11393 9267 11403 10151
rect 11011 6302 11403 9267
rect 11011 5994 11054 6302
rect 11362 5994 11403 6302
rect 3363 5573 3685 5842
rect 3363 5303 3391 5573
rect 1871 4831 2394 4841
rect 1871 4651 1916 4831
rect 2352 4651 2394 4831
rect 1871 4641 2394 4651
rect 357 2285 508 2307
rect 357 1109 364 2285
rect 500 1109 508 2285
rect 357 1087 508 1109
rect 856 913 1605 940
rect 856 891 884 913
rect 1576 891 1605 913
rect 856 755 882 891
rect 1578 755 1605 891
rect 856 733 884 755
rect 1576 733 1605 755
rect 856 706 1605 733
rect 2300 464 2394 4641
rect 2515 2703 3391 5303
rect 11011 5315 11403 5994
rect 11011 5007 11053 5315
rect 11361 5007 11403 5315
rect 2515 2459 2543 2703
rect 3363 2459 3391 2703
rect 2515 2403 3391 2459
rect 10573 1595 10732 4882
rect 11011 4451 11403 5007
rect 10976 4436 12119 4451
rect 10976 4064 11021 4436
rect 11393 4064 12119 4436
rect 10976 4050 12119 4064
rect 2484 1573 10732 1595
rect 2484 1457 2503 1573
rect 2683 1457 10732 1573
rect 2484 1436 10732 1457
rect 10952 2268 12119 2326
rect 2924 1256 3506 1305
rect 2924 756 2963 1256
rect 3463 803 3506 1256
rect 10952 803 11021 2268
rect 3463 756 11021 803
rect 2924 680 11021 756
rect 11393 1934 12119 2268
rect 11393 803 11921 1934
rect 11393 680 19235 803
rect 2924 578 19235 680
rect 11875 464 12216 483
rect 2300 452 12216 464
rect 2300 400 11891 452
rect 11943 400 11955 452
rect 12007 400 12019 452
rect 12071 400 12083 452
rect 12135 400 12147 452
rect 12199 400 12216 452
rect 2300 370 12216 400
rect 2478 238 3021 281
rect 2478 232 2534 238
rect 2970 232 3021 238
rect 2478 -64 2524 232
rect 2980 -64 3021 232
rect 2478 -70 2534 -64
rect 2970 -70 3021 -64
rect 2478 -114 3021 -70
rect 11278 238 11821 281
rect 11278 232 11334 238
rect 11770 232 11821 238
rect 11278 -64 11324 232
rect 11780 -64 11821 232
rect 11278 -70 11334 -64
rect 11770 -70 11821 -64
rect 11278 -114 11821 -70
<< via2 >>
rect 11058 10922 11354 11138
rect 364 1109 500 2285
rect 882 755 884 891
rect 884 755 1576 891
rect 1576 755 1578 891
rect 2524 -64 2534 232
rect 2534 -64 2970 232
rect 2970 -64 2980 232
rect 11324 -64 11334 232
rect 11334 -64 11770 232
rect 11770 -64 11780 232
<< metal3 >>
rect 11011 11142 11403 11182
rect 11011 10918 11054 11142
rect 11358 10918 11403 11142
rect 11011 10879 11403 10918
rect 337 2285 522 2321
rect 337 1109 364 2285
rect 500 1109 522 2285
rect 337 191 522 1109
rect 856 895 1605 940
rect 856 751 878 895
rect 1582 751 1605 895
rect 856 706 1605 751
rect 2478 236 3021 281
rect 2478 191 2520 236
rect 337 6 2520 191
rect 2478 -68 2520 6
rect 2984 -68 3021 236
rect 2478 -114 3021 -68
rect 11278 236 11821 281
rect 11278 -68 11320 236
rect 11784 -68 11821 236
rect 11278 -114 11821 -68
<< via3 >>
rect 11054 11138 11358 11142
rect 11054 10922 11058 11138
rect 11058 10922 11354 11138
rect 11354 10922 11358 11138
rect 11054 10918 11358 10922
rect 878 891 1582 895
rect 878 755 882 891
rect 882 755 1578 891
rect 1578 755 1582 891
rect 878 751 1582 755
rect 2520 232 2984 236
rect 2520 -64 2524 232
rect 2524 -64 2980 232
rect 2980 -64 2984 232
rect 2520 -68 2984 -64
rect 11320 232 11784 236
rect 11320 -64 11324 232
rect 11324 -64 11780 232
rect 11780 -64 11784 232
rect 11320 -68 11784 -64
<< metal4 >>
rect 0 11182 1039 11183
rect 0 10817 2236 11182
rect 11023 11142 11389 11170
rect 11023 10918 11054 11142
rect 11358 10918 11389 11142
rect 11023 10890 11389 10918
rect 0 10191 1606 10817
rect 857 895 1606 10191
rect 857 751 878 895
rect 1582 751 1606 895
rect 857 637 1606 751
rect 2478 236 3021 281
rect 2478 -68 2520 236
rect 2984 -68 3021 236
rect 2478 -114 3021 -68
rect 11278 236 11821 281
rect 11278 -68 11320 236
rect 11784 -68 11821 236
rect 11278 -114 11821 -68
<< via4 >>
rect 2634 -34 2870 202
rect 11434 -34 11670 202
<< metal5 >>
rect 2478 202 3021 281
rect 2478 -34 2634 202
rect 2870 -34 3021 202
rect 2478 -114 3021 -34
rect 11278 202 11871 281
rect 11278 -34 11434 202
rect 11670 -34 11871 202
rect 11278 -114 11871 -34
use hold_cap_array  hold_cap_array_0
timestamp 1699926577
transform 1 0 218 0 1 26439
box 1997 -26553 19047 -15257
use sky130_fd_pr__diode_pw2nd_05v5_L93GHW  sky130_fd_pr__diode_pw2nd_05v5_L93GHW_0
timestamp 1699926577
transform 1 0 778 0 1 9076
box -188 -188 188 188
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0
timestamp 1699926577
transform 0 1 409 -1 0 8738
box -66 -43 2178 1671
use balanced_switch  x1
timestamp 1699926577
transform -1 0 2730 0 1 2811
box 301 -2311 2543 1830
use follower_amp  x2
timestamp 1699926577
transform 1 0 8047 0 1 4397
box -4547 -3901 2817 6641
use follower_amp  x3
timestamp 1699926577
transform 1 0 16511 0 1 4407
box -4547 -3901 2817 6641
<< labels >>
flabel metal1 s 19269 4570 19469 4770 0 FreeSans 1 0 0 0 out
port 1 nsew
flabel metal1 s 0 5284 200 6015 0 FreeSans 1 0 0 0 vdd
port 2 nsew
flabel metal1 s 0 8901 200 9101 0 FreeSans 1 0 0 0 hold
port 3 nsew
flabel metal1 s 0 4986 200 5186 0 FreeSans 1 0 0 0 in
port 4 nsew
flabel metal4 s 0 10191 1039 11183 0 FreeSans 25 0 0 0 vss
port 5 nsew
flabel metal1 s 0 9612 804 9952 0 FreeSans 25 0 0 0 dvdd
port 6 nsew
flabel metal1 s 0 6152 788 6474 0 FreeSans 25 0 0 0 dvss
port 7 nsew
flabel metal1 s 0 4641 200 4841 0 FreeSans 1 0 0 0 ena
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 19469 11297
<< end >>
