magic
tech sky130A
magscale 1 2
timestamp 1699926577
<< pwell >>
rect -3349 -766 3349 766
<< mvnmos >>
rect -3131 318 -3031 518
rect -2973 318 -2873 518
rect -2815 318 -2715 518
rect -2657 318 -2557 518
rect -2499 318 -2399 518
rect -2341 318 -2241 518
rect -2183 318 -2083 518
rect -2025 318 -1925 518
rect -1867 318 -1767 518
rect -1709 318 -1609 518
rect -1551 318 -1451 518
rect -1393 318 -1293 518
rect -1235 318 -1135 518
rect -1077 318 -977 518
rect -919 318 -819 518
rect -761 318 -661 518
rect -603 318 -503 518
rect -445 318 -345 518
rect -287 318 -187 518
rect -129 318 -29 518
rect 29 318 129 518
rect 187 318 287 518
rect 345 318 445 518
rect 503 318 603 518
rect 661 318 761 518
rect 819 318 919 518
rect 977 318 1077 518
rect 1135 318 1235 518
rect 1293 318 1393 518
rect 1451 318 1551 518
rect 1609 318 1709 518
rect 1767 318 1867 518
rect 1925 318 2025 518
rect 2083 318 2183 518
rect 2241 318 2341 518
rect 2399 318 2499 518
rect 2557 318 2657 518
rect 2715 318 2815 518
rect 2873 318 2973 518
rect 3031 318 3131 518
rect -3131 -100 -3031 100
rect -2973 -100 -2873 100
rect -2815 -100 -2715 100
rect -2657 -100 -2557 100
rect -2499 -100 -2399 100
rect -2341 -100 -2241 100
rect -2183 -100 -2083 100
rect -2025 -100 -1925 100
rect -1867 -100 -1767 100
rect -1709 -100 -1609 100
rect -1551 -100 -1451 100
rect -1393 -100 -1293 100
rect -1235 -100 -1135 100
rect -1077 -100 -977 100
rect -919 -100 -819 100
rect -761 -100 -661 100
rect -603 -100 -503 100
rect -445 -100 -345 100
rect -287 -100 -187 100
rect -129 -100 -29 100
rect 29 -100 129 100
rect 187 -100 287 100
rect 345 -100 445 100
rect 503 -100 603 100
rect 661 -100 761 100
rect 819 -100 919 100
rect 977 -100 1077 100
rect 1135 -100 1235 100
rect 1293 -100 1393 100
rect 1451 -100 1551 100
rect 1609 -100 1709 100
rect 1767 -100 1867 100
rect 1925 -100 2025 100
rect 2083 -100 2183 100
rect 2241 -100 2341 100
rect 2399 -100 2499 100
rect 2557 -100 2657 100
rect 2715 -100 2815 100
rect 2873 -100 2973 100
rect 3031 -100 3131 100
rect -3131 -518 -3031 -318
rect -2973 -518 -2873 -318
rect -2815 -518 -2715 -318
rect -2657 -518 -2557 -318
rect -2499 -518 -2399 -318
rect -2341 -518 -2241 -318
rect -2183 -518 -2083 -318
rect -2025 -518 -1925 -318
rect -1867 -518 -1767 -318
rect -1709 -518 -1609 -318
rect -1551 -518 -1451 -318
rect -1393 -518 -1293 -318
rect -1235 -518 -1135 -318
rect -1077 -518 -977 -318
rect -919 -518 -819 -318
rect -761 -518 -661 -318
rect -603 -518 -503 -318
rect -445 -518 -345 -318
rect -287 -518 -187 -318
rect -129 -518 -29 -318
rect 29 -518 129 -318
rect 187 -518 287 -318
rect 345 -518 445 -318
rect 503 -518 603 -318
rect 661 -518 761 -318
rect 819 -518 919 -318
rect 977 -518 1077 -318
rect 1135 -518 1235 -318
rect 1293 -518 1393 -318
rect 1451 -518 1551 -318
rect 1609 -518 1709 -318
rect 1767 -518 1867 -318
rect 1925 -518 2025 -318
rect 2083 -518 2183 -318
rect 2241 -518 2341 -318
rect 2399 -518 2499 -318
rect 2557 -518 2657 -318
rect 2715 -518 2815 -318
rect 2873 -518 2973 -318
rect 3031 -518 3131 -318
<< mvndiff >>
rect -3189 503 -3131 518
rect -3189 469 -3177 503
rect -3143 469 -3131 503
rect -3189 435 -3131 469
rect -3189 401 -3177 435
rect -3143 401 -3131 435
rect -3189 367 -3131 401
rect -3189 333 -3177 367
rect -3143 333 -3131 367
rect -3189 318 -3131 333
rect -3031 503 -2973 518
rect -3031 469 -3019 503
rect -2985 469 -2973 503
rect -3031 435 -2973 469
rect -3031 401 -3019 435
rect -2985 401 -2973 435
rect -3031 367 -2973 401
rect -3031 333 -3019 367
rect -2985 333 -2973 367
rect -3031 318 -2973 333
rect -2873 503 -2815 518
rect -2873 469 -2861 503
rect -2827 469 -2815 503
rect -2873 435 -2815 469
rect -2873 401 -2861 435
rect -2827 401 -2815 435
rect -2873 367 -2815 401
rect -2873 333 -2861 367
rect -2827 333 -2815 367
rect -2873 318 -2815 333
rect -2715 503 -2657 518
rect -2715 469 -2703 503
rect -2669 469 -2657 503
rect -2715 435 -2657 469
rect -2715 401 -2703 435
rect -2669 401 -2657 435
rect -2715 367 -2657 401
rect -2715 333 -2703 367
rect -2669 333 -2657 367
rect -2715 318 -2657 333
rect -2557 503 -2499 518
rect -2557 469 -2545 503
rect -2511 469 -2499 503
rect -2557 435 -2499 469
rect -2557 401 -2545 435
rect -2511 401 -2499 435
rect -2557 367 -2499 401
rect -2557 333 -2545 367
rect -2511 333 -2499 367
rect -2557 318 -2499 333
rect -2399 503 -2341 518
rect -2399 469 -2387 503
rect -2353 469 -2341 503
rect -2399 435 -2341 469
rect -2399 401 -2387 435
rect -2353 401 -2341 435
rect -2399 367 -2341 401
rect -2399 333 -2387 367
rect -2353 333 -2341 367
rect -2399 318 -2341 333
rect -2241 503 -2183 518
rect -2241 469 -2229 503
rect -2195 469 -2183 503
rect -2241 435 -2183 469
rect -2241 401 -2229 435
rect -2195 401 -2183 435
rect -2241 367 -2183 401
rect -2241 333 -2229 367
rect -2195 333 -2183 367
rect -2241 318 -2183 333
rect -2083 503 -2025 518
rect -2083 469 -2071 503
rect -2037 469 -2025 503
rect -2083 435 -2025 469
rect -2083 401 -2071 435
rect -2037 401 -2025 435
rect -2083 367 -2025 401
rect -2083 333 -2071 367
rect -2037 333 -2025 367
rect -2083 318 -2025 333
rect -1925 503 -1867 518
rect -1925 469 -1913 503
rect -1879 469 -1867 503
rect -1925 435 -1867 469
rect -1925 401 -1913 435
rect -1879 401 -1867 435
rect -1925 367 -1867 401
rect -1925 333 -1913 367
rect -1879 333 -1867 367
rect -1925 318 -1867 333
rect -1767 503 -1709 518
rect -1767 469 -1755 503
rect -1721 469 -1709 503
rect -1767 435 -1709 469
rect -1767 401 -1755 435
rect -1721 401 -1709 435
rect -1767 367 -1709 401
rect -1767 333 -1755 367
rect -1721 333 -1709 367
rect -1767 318 -1709 333
rect -1609 503 -1551 518
rect -1609 469 -1597 503
rect -1563 469 -1551 503
rect -1609 435 -1551 469
rect -1609 401 -1597 435
rect -1563 401 -1551 435
rect -1609 367 -1551 401
rect -1609 333 -1597 367
rect -1563 333 -1551 367
rect -1609 318 -1551 333
rect -1451 503 -1393 518
rect -1451 469 -1439 503
rect -1405 469 -1393 503
rect -1451 435 -1393 469
rect -1451 401 -1439 435
rect -1405 401 -1393 435
rect -1451 367 -1393 401
rect -1451 333 -1439 367
rect -1405 333 -1393 367
rect -1451 318 -1393 333
rect -1293 503 -1235 518
rect -1293 469 -1281 503
rect -1247 469 -1235 503
rect -1293 435 -1235 469
rect -1293 401 -1281 435
rect -1247 401 -1235 435
rect -1293 367 -1235 401
rect -1293 333 -1281 367
rect -1247 333 -1235 367
rect -1293 318 -1235 333
rect -1135 503 -1077 518
rect -1135 469 -1123 503
rect -1089 469 -1077 503
rect -1135 435 -1077 469
rect -1135 401 -1123 435
rect -1089 401 -1077 435
rect -1135 367 -1077 401
rect -1135 333 -1123 367
rect -1089 333 -1077 367
rect -1135 318 -1077 333
rect -977 503 -919 518
rect -977 469 -965 503
rect -931 469 -919 503
rect -977 435 -919 469
rect -977 401 -965 435
rect -931 401 -919 435
rect -977 367 -919 401
rect -977 333 -965 367
rect -931 333 -919 367
rect -977 318 -919 333
rect -819 503 -761 518
rect -819 469 -807 503
rect -773 469 -761 503
rect -819 435 -761 469
rect -819 401 -807 435
rect -773 401 -761 435
rect -819 367 -761 401
rect -819 333 -807 367
rect -773 333 -761 367
rect -819 318 -761 333
rect -661 503 -603 518
rect -661 469 -649 503
rect -615 469 -603 503
rect -661 435 -603 469
rect -661 401 -649 435
rect -615 401 -603 435
rect -661 367 -603 401
rect -661 333 -649 367
rect -615 333 -603 367
rect -661 318 -603 333
rect -503 503 -445 518
rect -503 469 -491 503
rect -457 469 -445 503
rect -503 435 -445 469
rect -503 401 -491 435
rect -457 401 -445 435
rect -503 367 -445 401
rect -503 333 -491 367
rect -457 333 -445 367
rect -503 318 -445 333
rect -345 503 -287 518
rect -345 469 -333 503
rect -299 469 -287 503
rect -345 435 -287 469
rect -345 401 -333 435
rect -299 401 -287 435
rect -345 367 -287 401
rect -345 333 -333 367
rect -299 333 -287 367
rect -345 318 -287 333
rect -187 503 -129 518
rect -187 469 -175 503
rect -141 469 -129 503
rect -187 435 -129 469
rect -187 401 -175 435
rect -141 401 -129 435
rect -187 367 -129 401
rect -187 333 -175 367
rect -141 333 -129 367
rect -187 318 -129 333
rect -29 503 29 518
rect -29 469 -17 503
rect 17 469 29 503
rect -29 435 29 469
rect -29 401 -17 435
rect 17 401 29 435
rect -29 367 29 401
rect -29 333 -17 367
rect 17 333 29 367
rect -29 318 29 333
rect 129 503 187 518
rect 129 469 141 503
rect 175 469 187 503
rect 129 435 187 469
rect 129 401 141 435
rect 175 401 187 435
rect 129 367 187 401
rect 129 333 141 367
rect 175 333 187 367
rect 129 318 187 333
rect 287 503 345 518
rect 287 469 299 503
rect 333 469 345 503
rect 287 435 345 469
rect 287 401 299 435
rect 333 401 345 435
rect 287 367 345 401
rect 287 333 299 367
rect 333 333 345 367
rect 287 318 345 333
rect 445 503 503 518
rect 445 469 457 503
rect 491 469 503 503
rect 445 435 503 469
rect 445 401 457 435
rect 491 401 503 435
rect 445 367 503 401
rect 445 333 457 367
rect 491 333 503 367
rect 445 318 503 333
rect 603 503 661 518
rect 603 469 615 503
rect 649 469 661 503
rect 603 435 661 469
rect 603 401 615 435
rect 649 401 661 435
rect 603 367 661 401
rect 603 333 615 367
rect 649 333 661 367
rect 603 318 661 333
rect 761 503 819 518
rect 761 469 773 503
rect 807 469 819 503
rect 761 435 819 469
rect 761 401 773 435
rect 807 401 819 435
rect 761 367 819 401
rect 761 333 773 367
rect 807 333 819 367
rect 761 318 819 333
rect 919 503 977 518
rect 919 469 931 503
rect 965 469 977 503
rect 919 435 977 469
rect 919 401 931 435
rect 965 401 977 435
rect 919 367 977 401
rect 919 333 931 367
rect 965 333 977 367
rect 919 318 977 333
rect 1077 503 1135 518
rect 1077 469 1089 503
rect 1123 469 1135 503
rect 1077 435 1135 469
rect 1077 401 1089 435
rect 1123 401 1135 435
rect 1077 367 1135 401
rect 1077 333 1089 367
rect 1123 333 1135 367
rect 1077 318 1135 333
rect 1235 503 1293 518
rect 1235 469 1247 503
rect 1281 469 1293 503
rect 1235 435 1293 469
rect 1235 401 1247 435
rect 1281 401 1293 435
rect 1235 367 1293 401
rect 1235 333 1247 367
rect 1281 333 1293 367
rect 1235 318 1293 333
rect 1393 503 1451 518
rect 1393 469 1405 503
rect 1439 469 1451 503
rect 1393 435 1451 469
rect 1393 401 1405 435
rect 1439 401 1451 435
rect 1393 367 1451 401
rect 1393 333 1405 367
rect 1439 333 1451 367
rect 1393 318 1451 333
rect 1551 503 1609 518
rect 1551 469 1563 503
rect 1597 469 1609 503
rect 1551 435 1609 469
rect 1551 401 1563 435
rect 1597 401 1609 435
rect 1551 367 1609 401
rect 1551 333 1563 367
rect 1597 333 1609 367
rect 1551 318 1609 333
rect 1709 503 1767 518
rect 1709 469 1721 503
rect 1755 469 1767 503
rect 1709 435 1767 469
rect 1709 401 1721 435
rect 1755 401 1767 435
rect 1709 367 1767 401
rect 1709 333 1721 367
rect 1755 333 1767 367
rect 1709 318 1767 333
rect 1867 503 1925 518
rect 1867 469 1879 503
rect 1913 469 1925 503
rect 1867 435 1925 469
rect 1867 401 1879 435
rect 1913 401 1925 435
rect 1867 367 1925 401
rect 1867 333 1879 367
rect 1913 333 1925 367
rect 1867 318 1925 333
rect 2025 503 2083 518
rect 2025 469 2037 503
rect 2071 469 2083 503
rect 2025 435 2083 469
rect 2025 401 2037 435
rect 2071 401 2083 435
rect 2025 367 2083 401
rect 2025 333 2037 367
rect 2071 333 2083 367
rect 2025 318 2083 333
rect 2183 503 2241 518
rect 2183 469 2195 503
rect 2229 469 2241 503
rect 2183 435 2241 469
rect 2183 401 2195 435
rect 2229 401 2241 435
rect 2183 367 2241 401
rect 2183 333 2195 367
rect 2229 333 2241 367
rect 2183 318 2241 333
rect 2341 503 2399 518
rect 2341 469 2353 503
rect 2387 469 2399 503
rect 2341 435 2399 469
rect 2341 401 2353 435
rect 2387 401 2399 435
rect 2341 367 2399 401
rect 2341 333 2353 367
rect 2387 333 2399 367
rect 2341 318 2399 333
rect 2499 503 2557 518
rect 2499 469 2511 503
rect 2545 469 2557 503
rect 2499 435 2557 469
rect 2499 401 2511 435
rect 2545 401 2557 435
rect 2499 367 2557 401
rect 2499 333 2511 367
rect 2545 333 2557 367
rect 2499 318 2557 333
rect 2657 503 2715 518
rect 2657 469 2669 503
rect 2703 469 2715 503
rect 2657 435 2715 469
rect 2657 401 2669 435
rect 2703 401 2715 435
rect 2657 367 2715 401
rect 2657 333 2669 367
rect 2703 333 2715 367
rect 2657 318 2715 333
rect 2815 503 2873 518
rect 2815 469 2827 503
rect 2861 469 2873 503
rect 2815 435 2873 469
rect 2815 401 2827 435
rect 2861 401 2873 435
rect 2815 367 2873 401
rect 2815 333 2827 367
rect 2861 333 2873 367
rect 2815 318 2873 333
rect 2973 503 3031 518
rect 2973 469 2985 503
rect 3019 469 3031 503
rect 2973 435 3031 469
rect 2973 401 2985 435
rect 3019 401 3031 435
rect 2973 367 3031 401
rect 2973 333 2985 367
rect 3019 333 3031 367
rect 2973 318 3031 333
rect 3131 503 3189 518
rect 3131 469 3143 503
rect 3177 469 3189 503
rect 3131 435 3189 469
rect 3131 401 3143 435
rect 3177 401 3189 435
rect 3131 367 3189 401
rect 3131 333 3143 367
rect 3177 333 3189 367
rect 3131 318 3189 333
rect -3189 85 -3131 100
rect -3189 51 -3177 85
rect -3143 51 -3131 85
rect -3189 17 -3131 51
rect -3189 -17 -3177 17
rect -3143 -17 -3131 17
rect -3189 -51 -3131 -17
rect -3189 -85 -3177 -51
rect -3143 -85 -3131 -51
rect -3189 -100 -3131 -85
rect -3031 85 -2973 100
rect -3031 51 -3019 85
rect -2985 51 -2973 85
rect -3031 17 -2973 51
rect -3031 -17 -3019 17
rect -2985 -17 -2973 17
rect -3031 -51 -2973 -17
rect -3031 -85 -3019 -51
rect -2985 -85 -2973 -51
rect -3031 -100 -2973 -85
rect -2873 85 -2815 100
rect -2873 51 -2861 85
rect -2827 51 -2815 85
rect -2873 17 -2815 51
rect -2873 -17 -2861 17
rect -2827 -17 -2815 17
rect -2873 -51 -2815 -17
rect -2873 -85 -2861 -51
rect -2827 -85 -2815 -51
rect -2873 -100 -2815 -85
rect -2715 85 -2657 100
rect -2715 51 -2703 85
rect -2669 51 -2657 85
rect -2715 17 -2657 51
rect -2715 -17 -2703 17
rect -2669 -17 -2657 17
rect -2715 -51 -2657 -17
rect -2715 -85 -2703 -51
rect -2669 -85 -2657 -51
rect -2715 -100 -2657 -85
rect -2557 85 -2499 100
rect -2557 51 -2545 85
rect -2511 51 -2499 85
rect -2557 17 -2499 51
rect -2557 -17 -2545 17
rect -2511 -17 -2499 17
rect -2557 -51 -2499 -17
rect -2557 -85 -2545 -51
rect -2511 -85 -2499 -51
rect -2557 -100 -2499 -85
rect -2399 85 -2341 100
rect -2399 51 -2387 85
rect -2353 51 -2341 85
rect -2399 17 -2341 51
rect -2399 -17 -2387 17
rect -2353 -17 -2341 17
rect -2399 -51 -2341 -17
rect -2399 -85 -2387 -51
rect -2353 -85 -2341 -51
rect -2399 -100 -2341 -85
rect -2241 85 -2183 100
rect -2241 51 -2229 85
rect -2195 51 -2183 85
rect -2241 17 -2183 51
rect -2241 -17 -2229 17
rect -2195 -17 -2183 17
rect -2241 -51 -2183 -17
rect -2241 -85 -2229 -51
rect -2195 -85 -2183 -51
rect -2241 -100 -2183 -85
rect -2083 85 -2025 100
rect -2083 51 -2071 85
rect -2037 51 -2025 85
rect -2083 17 -2025 51
rect -2083 -17 -2071 17
rect -2037 -17 -2025 17
rect -2083 -51 -2025 -17
rect -2083 -85 -2071 -51
rect -2037 -85 -2025 -51
rect -2083 -100 -2025 -85
rect -1925 85 -1867 100
rect -1925 51 -1913 85
rect -1879 51 -1867 85
rect -1925 17 -1867 51
rect -1925 -17 -1913 17
rect -1879 -17 -1867 17
rect -1925 -51 -1867 -17
rect -1925 -85 -1913 -51
rect -1879 -85 -1867 -51
rect -1925 -100 -1867 -85
rect -1767 85 -1709 100
rect -1767 51 -1755 85
rect -1721 51 -1709 85
rect -1767 17 -1709 51
rect -1767 -17 -1755 17
rect -1721 -17 -1709 17
rect -1767 -51 -1709 -17
rect -1767 -85 -1755 -51
rect -1721 -85 -1709 -51
rect -1767 -100 -1709 -85
rect -1609 85 -1551 100
rect -1609 51 -1597 85
rect -1563 51 -1551 85
rect -1609 17 -1551 51
rect -1609 -17 -1597 17
rect -1563 -17 -1551 17
rect -1609 -51 -1551 -17
rect -1609 -85 -1597 -51
rect -1563 -85 -1551 -51
rect -1609 -100 -1551 -85
rect -1451 85 -1393 100
rect -1451 51 -1439 85
rect -1405 51 -1393 85
rect -1451 17 -1393 51
rect -1451 -17 -1439 17
rect -1405 -17 -1393 17
rect -1451 -51 -1393 -17
rect -1451 -85 -1439 -51
rect -1405 -85 -1393 -51
rect -1451 -100 -1393 -85
rect -1293 85 -1235 100
rect -1293 51 -1281 85
rect -1247 51 -1235 85
rect -1293 17 -1235 51
rect -1293 -17 -1281 17
rect -1247 -17 -1235 17
rect -1293 -51 -1235 -17
rect -1293 -85 -1281 -51
rect -1247 -85 -1235 -51
rect -1293 -100 -1235 -85
rect -1135 85 -1077 100
rect -1135 51 -1123 85
rect -1089 51 -1077 85
rect -1135 17 -1077 51
rect -1135 -17 -1123 17
rect -1089 -17 -1077 17
rect -1135 -51 -1077 -17
rect -1135 -85 -1123 -51
rect -1089 -85 -1077 -51
rect -1135 -100 -1077 -85
rect -977 85 -919 100
rect -977 51 -965 85
rect -931 51 -919 85
rect -977 17 -919 51
rect -977 -17 -965 17
rect -931 -17 -919 17
rect -977 -51 -919 -17
rect -977 -85 -965 -51
rect -931 -85 -919 -51
rect -977 -100 -919 -85
rect -819 85 -761 100
rect -819 51 -807 85
rect -773 51 -761 85
rect -819 17 -761 51
rect -819 -17 -807 17
rect -773 -17 -761 17
rect -819 -51 -761 -17
rect -819 -85 -807 -51
rect -773 -85 -761 -51
rect -819 -100 -761 -85
rect -661 85 -603 100
rect -661 51 -649 85
rect -615 51 -603 85
rect -661 17 -603 51
rect -661 -17 -649 17
rect -615 -17 -603 17
rect -661 -51 -603 -17
rect -661 -85 -649 -51
rect -615 -85 -603 -51
rect -661 -100 -603 -85
rect -503 85 -445 100
rect -503 51 -491 85
rect -457 51 -445 85
rect -503 17 -445 51
rect -503 -17 -491 17
rect -457 -17 -445 17
rect -503 -51 -445 -17
rect -503 -85 -491 -51
rect -457 -85 -445 -51
rect -503 -100 -445 -85
rect -345 85 -287 100
rect -345 51 -333 85
rect -299 51 -287 85
rect -345 17 -287 51
rect -345 -17 -333 17
rect -299 -17 -287 17
rect -345 -51 -287 -17
rect -345 -85 -333 -51
rect -299 -85 -287 -51
rect -345 -100 -287 -85
rect -187 85 -129 100
rect -187 51 -175 85
rect -141 51 -129 85
rect -187 17 -129 51
rect -187 -17 -175 17
rect -141 -17 -129 17
rect -187 -51 -129 -17
rect -187 -85 -175 -51
rect -141 -85 -129 -51
rect -187 -100 -129 -85
rect -29 85 29 100
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -100 29 -85
rect 129 85 187 100
rect 129 51 141 85
rect 175 51 187 85
rect 129 17 187 51
rect 129 -17 141 17
rect 175 -17 187 17
rect 129 -51 187 -17
rect 129 -85 141 -51
rect 175 -85 187 -51
rect 129 -100 187 -85
rect 287 85 345 100
rect 287 51 299 85
rect 333 51 345 85
rect 287 17 345 51
rect 287 -17 299 17
rect 333 -17 345 17
rect 287 -51 345 -17
rect 287 -85 299 -51
rect 333 -85 345 -51
rect 287 -100 345 -85
rect 445 85 503 100
rect 445 51 457 85
rect 491 51 503 85
rect 445 17 503 51
rect 445 -17 457 17
rect 491 -17 503 17
rect 445 -51 503 -17
rect 445 -85 457 -51
rect 491 -85 503 -51
rect 445 -100 503 -85
rect 603 85 661 100
rect 603 51 615 85
rect 649 51 661 85
rect 603 17 661 51
rect 603 -17 615 17
rect 649 -17 661 17
rect 603 -51 661 -17
rect 603 -85 615 -51
rect 649 -85 661 -51
rect 603 -100 661 -85
rect 761 85 819 100
rect 761 51 773 85
rect 807 51 819 85
rect 761 17 819 51
rect 761 -17 773 17
rect 807 -17 819 17
rect 761 -51 819 -17
rect 761 -85 773 -51
rect 807 -85 819 -51
rect 761 -100 819 -85
rect 919 85 977 100
rect 919 51 931 85
rect 965 51 977 85
rect 919 17 977 51
rect 919 -17 931 17
rect 965 -17 977 17
rect 919 -51 977 -17
rect 919 -85 931 -51
rect 965 -85 977 -51
rect 919 -100 977 -85
rect 1077 85 1135 100
rect 1077 51 1089 85
rect 1123 51 1135 85
rect 1077 17 1135 51
rect 1077 -17 1089 17
rect 1123 -17 1135 17
rect 1077 -51 1135 -17
rect 1077 -85 1089 -51
rect 1123 -85 1135 -51
rect 1077 -100 1135 -85
rect 1235 85 1293 100
rect 1235 51 1247 85
rect 1281 51 1293 85
rect 1235 17 1293 51
rect 1235 -17 1247 17
rect 1281 -17 1293 17
rect 1235 -51 1293 -17
rect 1235 -85 1247 -51
rect 1281 -85 1293 -51
rect 1235 -100 1293 -85
rect 1393 85 1451 100
rect 1393 51 1405 85
rect 1439 51 1451 85
rect 1393 17 1451 51
rect 1393 -17 1405 17
rect 1439 -17 1451 17
rect 1393 -51 1451 -17
rect 1393 -85 1405 -51
rect 1439 -85 1451 -51
rect 1393 -100 1451 -85
rect 1551 85 1609 100
rect 1551 51 1563 85
rect 1597 51 1609 85
rect 1551 17 1609 51
rect 1551 -17 1563 17
rect 1597 -17 1609 17
rect 1551 -51 1609 -17
rect 1551 -85 1563 -51
rect 1597 -85 1609 -51
rect 1551 -100 1609 -85
rect 1709 85 1767 100
rect 1709 51 1721 85
rect 1755 51 1767 85
rect 1709 17 1767 51
rect 1709 -17 1721 17
rect 1755 -17 1767 17
rect 1709 -51 1767 -17
rect 1709 -85 1721 -51
rect 1755 -85 1767 -51
rect 1709 -100 1767 -85
rect 1867 85 1925 100
rect 1867 51 1879 85
rect 1913 51 1925 85
rect 1867 17 1925 51
rect 1867 -17 1879 17
rect 1913 -17 1925 17
rect 1867 -51 1925 -17
rect 1867 -85 1879 -51
rect 1913 -85 1925 -51
rect 1867 -100 1925 -85
rect 2025 85 2083 100
rect 2025 51 2037 85
rect 2071 51 2083 85
rect 2025 17 2083 51
rect 2025 -17 2037 17
rect 2071 -17 2083 17
rect 2025 -51 2083 -17
rect 2025 -85 2037 -51
rect 2071 -85 2083 -51
rect 2025 -100 2083 -85
rect 2183 85 2241 100
rect 2183 51 2195 85
rect 2229 51 2241 85
rect 2183 17 2241 51
rect 2183 -17 2195 17
rect 2229 -17 2241 17
rect 2183 -51 2241 -17
rect 2183 -85 2195 -51
rect 2229 -85 2241 -51
rect 2183 -100 2241 -85
rect 2341 85 2399 100
rect 2341 51 2353 85
rect 2387 51 2399 85
rect 2341 17 2399 51
rect 2341 -17 2353 17
rect 2387 -17 2399 17
rect 2341 -51 2399 -17
rect 2341 -85 2353 -51
rect 2387 -85 2399 -51
rect 2341 -100 2399 -85
rect 2499 85 2557 100
rect 2499 51 2511 85
rect 2545 51 2557 85
rect 2499 17 2557 51
rect 2499 -17 2511 17
rect 2545 -17 2557 17
rect 2499 -51 2557 -17
rect 2499 -85 2511 -51
rect 2545 -85 2557 -51
rect 2499 -100 2557 -85
rect 2657 85 2715 100
rect 2657 51 2669 85
rect 2703 51 2715 85
rect 2657 17 2715 51
rect 2657 -17 2669 17
rect 2703 -17 2715 17
rect 2657 -51 2715 -17
rect 2657 -85 2669 -51
rect 2703 -85 2715 -51
rect 2657 -100 2715 -85
rect 2815 85 2873 100
rect 2815 51 2827 85
rect 2861 51 2873 85
rect 2815 17 2873 51
rect 2815 -17 2827 17
rect 2861 -17 2873 17
rect 2815 -51 2873 -17
rect 2815 -85 2827 -51
rect 2861 -85 2873 -51
rect 2815 -100 2873 -85
rect 2973 85 3031 100
rect 2973 51 2985 85
rect 3019 51 3031 85
rect 2973 17 3031 51
rect 2973 -17 2985 17
rect 3019 -17 3031 17
rect 2973 -51 3031 -17
rect 2973 -85 2985 -51
rect 3019 -85 3031 -51
rect 2973 -100 3031 -85
rect 3131 85 3189 100
rect 3131 51 3143 85
rect 3177 51 3189 85
rect 3131 17 3189 51
rect 3131 -17 3143 17
rect 3177 -17 3189 17
rect 3131 -51 3189 -17
rect 3131 -85 3143 -51
rect 3177 -85 3189 -51
rect 3131 -100 3189 -85
rect -3189 -333 -3131 -318
rect -3189 -367 -3177 -333
rect -3143 -367 -3131 -333
rect -3189 -401 -3131 -367
rect -3189 -435 -3177 -401
rect -3143 -435 -3131 -401
rect -3189 -469 -3131 -435
rect -3189 -503 -3177 -469
rect -3143 -503 -3131 -469
rect -3189 -518 -3131 -503
rect -3031 -333 -2973 -318
rect -3031 -367 -3019 -333
rect -2985 -367 -2973 -333
rect -3031 -401 -2973 -367
rect -3031 -435 -3019 -401
rect -2985 -435 -2973 -401
rect -3031 -469 -2973 -435
rect -3031 -503 -3019 -469
rect -2985 -503 -2973 -469
rect -3031 -518 -2973 -503
rect -2873 -333 -2815 -318
rect -2873 -367 -2861 -333
rect -2827 -367 -2815 -333
rect -2873 -401 -2815 -367
rect -2873 -435 -2861 -401
rect -2827 -435 -2815 -401
rect -2873 -469 -2815 -435
rect -2873 -503 -2861 -469
rect -2827 -503 -2815 -469
rect -2873 -518 -2815 -503
rect -2715 -333 -2657 -318
rect -2715 -367 -2703 -333
rect -2669 -367 -2657 -333
rect -2715 -401 -2657 -367
rect -2715 -435 -2703 -401
rect -2669 -435 -2657 -401
rect -2715 -469 -2657 -435
rect -2715 -503 -2703 -469
rect -2669 -503 -2657 -469
rect -2715 -518 -2657 -503
rect -2557 -333 -2499 -318
rect -2557 -367 -2545 -333
rect -2511 -367 -2499 -333
rect -2557 -401 -2499 -367
rect -2557 -435 -2545 -401
rect -2511 -435 -2499 -401
rect -2557 -469 -2499 -435
rect -2557 -503 -2545 -469
rect -2511 -503 -2499 -469
rect -2557 -518 -2499 -503
rect -2399 -333 -2341 -318
rect -2399 -367 -2387 -333
rect -2353 -367 -2341 -333
rect -2399 -401 -2341 -367
rect -2399 -435 -2387 -401
rect -2353 -435 -2341 -401
rect -2399 -469 -2341 -435
rect -2399 -503 -2387 -469
rect -2353 -503 -2341 -469
rect -2399 -518 -2341 -503
rect -2241 -333 -2183 -318
rect -2241 -367 -2229 -333
rect -2195 -367 -2183 -333
rect -2241 -401 -2183 -367
rect -2241 -435 -2229 -401
rect -2195 -435 -2183 -401
rect -2241 -469 -2183 -435
rect -2241 -503 -2229 -469
rect -2195 -503 -2183 -469
rect -2241 -518 -2183 -503
rect -2083 -333 -2025 -318
rect -2083 -367 -2071 -333
rect -2037 -367 -2025 -333
rect -2083 -401 -2025 -367
rect -2083 -435 -2071 -401
rect -2037 -435 -2025 -401
rect -2083 -469 -2025 -435
rect -2083 -503 -2071 -469
rect -2037 -503 -2025 -469
rect -2083 -518 -2025 -503
rect -1925 -333 -1867 -318
rect -1925 -367 -1913 -333
rect -1879 -367 -1867 -333
rect -1925 -401 -1867 -367
rect -1925 -435 -1913 -401
rect -1879 -435 -1867 -401
rect -1925 -469 -1867 -435
rect -1925 -503 -1913 -469
rect -1879 -503 -1867 -469
rect -1925 -518 -1867 -503
rect -1767 -333 -1709 -318
rect -1767 -367 -1755 -333
rect -1721 -367 -1709 -333
rect -1767 -401 -1709 -367
rect -1767 -435 -1755 -401
rect -1721 -435 -1709 -401
rect -1767 -469 -1709 -435
rect -1767 -503 -1755 -469
rect -1721 -503 -1709 -469
rect -1767 -518 -1709 -503
rect -1609 -333 -1551 -318
rect -1609 -367 -1597 -333
rect -1563 -367 -1551 -333
rect -1609 -401 -1551 -367
rect -1609 -435 -1597 -401
rect -1563 -435 -1551 -401
rect -1609 -469 -1551 -435
rect -1609 -503 -1597 -469
rect -1563 -503 -1551 -469
rect -1609 -518 -1551 -503
rect -1451 -333 -1393 -318
rect -1451 -367 -1439 -333
rect -1405 -367 -1393 -333
rect -1451 -401 -1393 -367
rect -1451 -435 -1439 -401
rect -1405 -435 -1393 -401
rect -1451 -469 -1393 -435
rect -1451 -503 -1439 -469
rect -1405 -503 -1393 -469
rect -1451 -518 -1393 -503
rect -1293 -333 -1235 -318
rect -1293 -367 -1281 -333
rect -1247 -367 -1235 -333
rect -1293 -401 -1235 -367
rect -1293 -435 -1281 -401
rect -1247 -435 -1235 -401
rect -1293 -469 -1235 -435
rect -1293 -503 -1281 -469
rect -1247 -503 -1235 -469
rect -1293 -518 -1235 -503
rect -1135 -333 -1077 -318
rect -1135 -367 -1123 -333
rect -1089 -367 -1077 -333
rect -1135 -401 -1077 -367
rect -1135 -435 -1123 -401
rect -1089 -435 -1077 -401
rect -1135 -469 -1077 -435
rect -1135 -503 -1123 -469
rect -1089 -503 -1077 -469
rect -1135 -518 -1077 -503
rect -977 -333 -919 -318
rect -977 -367 -965 -333
rect -931 -367 -919 -333
rect -977 -401 -919 -367
rect -977 -435 -965 -401
rect -931 -435 -919 -401
rect -977 -469 -919 -435
rect -977 -503 -965 -469
rect -931 -503 -919 -469
rect -977 -518 -919 -503
rect -819 -333 -761 -318
rect -819 -367 -807 -333
rect -773 -367 -761 -333
rect -819 -401 -761 -367
rect -819 -435 -807 -401
rect -773 -435 -761 -401
rect -819 -469 -761 -435
rect -819 -503 -807 -469
rect -773 -503 -761 -469
rect -819 -518 -761 -503
rect -661 -333 -603 -318
rect -661 -367 -649 -333
rect -615 -367 -603 -333
rect -661 -401 -603 -367
rect -661 -435 -649 -401
rect -615 -435 -603 -401
rect -661 -469 -603 -435
rect -661 -503 -649 -469
rect -615 -503 -603 -469
rect -661 -518 -603 -503
rect -503 -333 -445 -318
rect -503 -367 -491 -333
rect -457 -367 -445 -333
rect -503 -401 -445 -367
rect -503 -435 -491 -401
rect -457 -435 -445 -401
rect -503 -469 -445 -435
rect -503 -503 -491 -469
rect -457 -503 -445 -469
rect -503 -518 -445 -503
rect -345 -333 -287 -318
rect -345 -367 -333 -333
rect -299 -367 -287 -333
rect -345 -401 -287 -367
rect -345 -435 -333 -401
rect -299 -435 -287 -401
rect -345 -469 -287 -435
rect -345 -503 -333 -469
rect -299 -503 -287 -469
rect -345 -518 -287 -503
rect -187 -333 -129 -318
rect -187 -367 -175 -333
rect -141 -367 -129 -333
rect -187 -401 -129 -367
rect -187 -435 -175 -401
rect -141 -435 -129 -401
rect -187 -469 -129 -435
rect -187 -503 -175 -469
rect -141 -503 -129 -469
rect -187 -518 -129 -503
rect -29 -333 29 -318
rect -29 -367 -17 -333
rect 17 -367 29 -333
rect -29 -401 29 -367
rect -29 -435 -17 -401
rect 17 -435 29 -401
rect -29 -469 29 -435
rect -29 -503 -17 -469
rect 17 -503 29 -469
rect -29 -518 29 -503
rect 129 -333 187 -318
rect 129 -367 141 -333
rect 175 -367 187 -333
rect 129 -401 187 -367
rect 129 -435 141 -401
rect 175 -435 187 -401
rect 129 -469 187 -435
rect 129 -503 141 -469
rect 175 -503 187 -469
rect 129 -518 187 -503
rect 287 -333 345 -318
rect 287 -367 299 -333
rect 333 -367 345 -333
rect 287 -401 345 -367
rect 287 -435 299 -401
rect 333 -435 345 -401
rect 287 -469 345 -435
rect 287 -503 299 -469
rect 333 -503 345 -469
rect 287 -518 345 -503
rect 445 -333 503 -318
rect 445 -367 457 -333
rect 491 -367 503 -333
rect 445 -401 503 -367
rect 445 -435 457 -401
rect 491 -435 503 -401
rect 445 -469 503 -435
rect 445 -503 457 -469
rect 491 -503 503 -469
rect 445 -518 503 -503
rect 603 -333 661 -318
rect 603 -367 615 -333
rect 649 -367 661 -333
rect 603 -401 661 -367
rect 603 -435 615 -401
rect 649 -435 661 -401
rect 603 -469 661 -435
rect 603 -503 615 -469
rect 649 -503 661 -469
rect 603 -518 661 -503
rect 761 -333 819 -318
rect 761 -367 773 -333
rect 807 -367 819 -333
rect 761 -401 819 -367
rect 761 -435 773 -401
rect 807 -435 819 -401
rect 761 -469 819 -435
rect 761 -503 773 -469
rect 807 -503 819 -469
rect 761 -518 819 -503
rect 919 -333 977 -318
rect 919 -367 931 -333
rect 965 -367 977 -333
rect 919 -401 977 -367
rect 919 -435 931 -401
rect 965 -435 977 -401
rect 919 -469 977 -435
rect 919 -503 931 -469
rect 965 -503 977 -469
rect 919 -518 977 -503
rect 1077 -333 1135 -318
rect 1077 -367 1089 -333
rect 1123 -367 1135 -333
rect 1077 -401 1135 -367
rect 1077 -435 1089 -401
rect 1123 -435 1135 -401
rect 1077 -469 1135 -435
rect 1077 -503 1089 -469
rect 1123 -503 1135 -469
rect 1077 -518 1135 -503
rect 1235 -333 1293 -318
rect 1235 -367 1247 -333
rect 1281 -367 1293 -333
rect 1235 -401 1293 -367
rect 1235 -435 1247 -401
rect 1281 -435 1293 -401
rect 1235 -469 1293 -435
rect 1235 -503 1247 -469
rect 1281 -503 1293 -469
rect 1235 -518 1293 -503
rect 1393 -333 1451 -318
rect 1393 -367 1405 -333
rect 1439 -367 1451 -333
rect 1393 -401 1451 -367
rect 1393 -435 1405 -401
rect 1439 -435 1451 -401
rect 1393 -469 1451 -435
rect 1393 -503 1405 -469
rect 1439 -503 1451 -469
rect 1393 -518 1451 -503
rect 1551 -333 1609 -318
rect 1551 -367 1563 -333
rect 1597 -367 1609 -333
rect 1551 -401 1609 -367
rect 1551 -435 1563 -401
rect 1597 -435 1609 -401
rect 1551 -469 1609 -435
rect 1551 -503 1563 -469
rect 1597 -503 1609 -469
rect 1551 -518 1609 -503
rect 1709 -333 1767 -318
rect 1709 -367 1721 -333
rect 1755 -367 1767 -333
rect 1709 -401 1767 -367
rect 1709 -435 1721 -401
rect 1755 -435 1767 -401
rect 1709 -469 1767 -435
rect 1709 -503 1721 -469
rect 1755 -503 1767 -469
rect 1709 -518 1767 -503
rect 1867 -333 1925 -318
rect 1867 -367 1879 -333
rect 1913 -367 1925 -333
rect 1867 -401 1925 -367
rect 1867 -435 1879 -401
rect 1913 -435 1925 -401
rect 1867 -469 1925 -435
rect 1867 -503 1879 -469
rect 1913 -503 1925 -469
rect 1867 -518 1925 -503
rect 2025 -333 2083 -318
rect 2025 -367 2037 -333
rect 2071 -367 2083 -333
rect 2025 -401 2083 -367
rect 2025 -435 2037 -401
rect 2071 -435 2083 -401
rect 2025 -469 2083 -435
rect 2025 -503 2037 -469
rect 2071 -503 2083 -469
rect 2025 -518 2083 -503
rect 2183 -333 2241 -318
rect 2183 -367 2195 -333
rect 2229 -367 2241 -333
rect 2183 -401 2241 -367
rect 2183 -435 2195 -401
rect 2229 -435 2241 -401
rect 2183 -469 2241 -435
rect 2183 -503 2195 -469
rect 2229 -503 2241 -469
rect 2183 -518 2241 -503
rect 2341 -333 2399 -318
rect 2341 -367 2353 -333
rect 2387 -367 2399 -333
rect 2341 -401 2399 -367
rect 2341 -435 2353 -401
rect 2387 -435 2399 -401
rect 2341 -469 2399 -435
rect 2341 -503 2353 -469
rect 2387 -503 2399 -469
rect 2341 -518 2399 -503
rect 2499 -333 2557 -318
rect 2499 -367 2511 -333
rect 2545 -367 2557 -333
rect 2499 -401 2557 -367
rect 2499 -435 2511 -401
rect 2545 -435 2557 -401
rect 2499 -469 2557 -435
rect 2499 -503 2511 -469
rect 2545 -503 2557 -469
rect 2499 -518 2557 -503
rect 2657 -333 2715 -318
rect 2657 -367 2669 -333
rect 2703 -367 2715 -333
rect 2657 -401 2715 -367
rect 2657 -435 2669 -401
rect 2703 -435 2715 -401
rect 2657 -469 2715 -435
rect 2657 -503 2669 -469
rect 2703 -503 2715 -469
rect 2657 -518 2715 -503
rect 2815 -333 2873 -318
rect 2815 -367 2827 -333
rect 2861 -367 2873 -333
rect 2815 -401 2873 -367
rect 2815 -435 2827 -401
rect 2861 -435 2873 -401
rect 2815 -469 2873 -435
rect 2815 -503 2827 -469
rect 2861 -503 2873 -469
rect 2815 -518 2873 -503
rect 2973 -333 3031 -318
rect 2973 -367 2985 -333
rect 3019 -367 3031 -333
rect 2973 -401 3031 -367
rect 2973 -435 2985 -401
rect 3019 -435 3031 -401
rect 2973 -469 3031 -435
rect 2973 -503 2985 -469
rect 3019 -503 3031 -469
rect 2973 -518 3031 -503
rect 3131 -333 3189 -318
rect 3131 -367 3143 -333
rect 3177 -367 3189 -333
rect 3131 -401 3189 -367
rect 3131 -435 3143 -401
rect 3177 -435 3189 -401
rect 3131 -469 3189 -435
rect 3131 -503 3143 -469
rect 3177 -503 3189 -469
rect 3131 -518 3189 -503
<< mvndiffc >>
rect -3177 469 -3143 503
rect -3177 401 -3143 435
rect -3177 333 -3143 367
rect -3019 469 -2985 503
rect -3019 401 -2985 435
rect -3019 333 -2985 367
rect -2861 469 -2827 503
rect -2861 401 -2827 435
rect -2861 333 -2827 367
rect -2703 469 -2669 503
rect -2703 401 -2669 435
rect -2703 333 -2669 367
rect -2545 469 -2511 503
rect -2545 401 -2511 435
rect -2545 333 -2511 367
rect -2387 469 -2353 503
rect -2387 401 -2353 435
rect -2387 333 -2353 367
rect -2229 469 -2195 503
rect -2229 401 -2195 435
rect -2229 333 -2195 367
rect -2071 469 -2037 503
rect -2071 401 -2037 435
rect -2071 333 -2037 367
rect -1913 469 -1879 503
rect -1913 401 -1879 435
rect -1913 333 -1879 367
rect -1755 469 -1721 503
rect -1755 401 -1721 435
rect -1755 333 -1721 367
rect -1597 469 -1563 503
rect -1597 401 -1563 435
rect -1597 333 -1563 367
rect -1439 469 -1405 503
rect -1439 401 -1405 435
rect -1439 333 -1405 367
rect -1281 469 -1247 503
rect -1281 401 -1247 435
rect -1281 333 -1247 367
rect -1123 469 -1089 503
rect -1123 401 -1089 435
rect -1123 333 -1089 367
rect -965 469 -931 503
rect -965 401 -931 435
rect -965 333 -931 367
rect -807 469 -773 503
rect -807 401 -773 435
rect -807 333 -773 367
rect -649 469 -615 503
rect -649 401 -615 435
rect -649 333 -615 367
rect -491 469 -457 503
rect -491 401 -457 435
rect -491 333 -457 367
rect -333 469 -299 503
rect -333 401 -299 435
rect -333 333 -299 367
rect -175 469 -141 503
rect -175 401 -141 435
rect -175 333 -141 367
rect -17 469 17 503
rect -17 401 17 435
rect -17 333 17 367
rect 141 469 175 503
rect 141 401 175 435
rect 141 333 175 367
rect 299 469 333 503
rect 299 401 333 435
rect 299 333 333 367
rect 457 469 491 503
rect 457 401 491 435
rect 457 333 491 367
rect 615 469 649 503
rect 615 401 649 435
rect 615 333 649 367
rect 773 469 807 503
rect 773 401 807 435
rect 773 333 807 367
rect 931 469 965 503
rect 931 401 965 435
rect 931 333 965 367
rect 1089 469 1123 503
rect 1089 401 1123 435
rect 1089 333 1123 367
rect 1247 469 1281 503
rect 1247 401 1281 435
rect 1247 333 1281 367
rect 1405 469 1439 503
rect 1405 401 1439 435
rect 1405 333 1439 367
rect 1563 469 1597 503
rect 1563 401 1597 435
rect 1563 333 1597 367
rect 1721 469 1755 503
rect 1721 401 1755 435
rect 1721 333 1755 367
rect 1879 469 1913 503
rect 1879 401 1913 435
rect 1879 333 1913 367
rect 2037 469 2071 503
rect 2037 401 2071 435
rect 2037 333 2071 367
rect 2195 469 2229 503
rect 2195 401 2229 435
rect 2195 333 2229 367
rect 2353 469 2387 503
rect 2353 401 2387 435
rect 2353 333 2387 367
rect 2511 469 2545 503
rect 2511 401 2545 435
rect 2511 333 2545 367
rect 2669 469 2703 503
rect 2669 401 2703 435
rect 2669 333 2703 367
rect 2827 469 2861 503
rect 2827 401 2861 435
rect 2827 333 2861 367
rect 2985 469 3019 503
rect 2985 401 3019 435
rect 2985 333 3019 367
rect 3143 469 3177 503
rect 3143 401 3177 435
rect 3143 333 3177 367
rect -3177 51 -3143 85
rect -3177 -17 -3143 17
rect -3177 -85 -3143 -51
rect -3019 51 -2985 85
rect -3019 -17 -2985 17
rect -3019 -85 -2985 -51
rect -2861 51 -2827 85
rect -2861 -17 -2827 17
rect -2861 -85 -2827 -51
rect -2703 51 -2669 85
rect -2703 -17 -2669 17
rect -2703 -85 -2669 -51
rect -2545 51 -2511 85
rect -2545 -17 -2511 17
rect -2545 -85 -2511 -51
rect -2387 51 -2353 85
rect -2387 -17 -2353 17
rect -2387 -85 -2353 -51
rect -2229 51 -2195 85
rect -2229 -17 -2195 17
rect -2229 -85 -2195 -51
rect -2071 51 -2037 85
rect -2071 -17 -2037 17
rect -2071 -85 -2037 -51
rect -1913 51 -1879 85
rect -1913 -17 -1879 17
rect -1913 -85 -1879 -51
rect -1755 51 -1721 85
rect -1755 -17 -1721 17
rect -1755 -85 -1721 -51
rect -1597 51 -1563 85
rect -1597 -17 -1563 17
rect -1597 -85 -1563 -51
rect -1439 51 -1405 85
rect -1439 -17 -1405 17
rect -1439 -85 -1405 -51
rect -1281 51 -1247 85
rect -1281 -17 -1247 17
rect -1281 -85 -1247 -51
rect -1123 51 -1089 85
rect -1123 -17 -1089 17
rect -1123 -85 -1089 -51
rect -965 51 -931 85
rect -965 -17 -931 17
rect -965 -85 -931 -51
rect -807 51 -773 85
rect -807 -17 -773 17
rect -807 -85 -773 -51
rect -649 51 -615 85
rect -649 -17 -615 17
rect -649 -85 -615 -51
rect -491 51 -457 85
rect -491 -17 -457 17
rect -491 -85 -457 -51
rect -333 51 -299 85
rect -333 -17 -299 17
rect -333 -85 -299 -51
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect 299 51 333 85
rect 299 -17 333 17
rect 299 -85 333 -51
rect 457 51 491 85
rect 457 -17 491 17
rect 457 -85 491 -51
rect 615 51 649 85
rect 615 -17 649 17
rect 615 -85 649 -51
rect 773 51 807 85
rect 773 -17 807 17
rect 773 -85 807 -51
rect 931 51 965 85
rect 931 -17 965 17
rect 931 -85 965 -51
rect 1089 51 1123 85
rect 1089 -17 1123 17
rect 1089 -85 1123 -51
rect 1247 51 1281 85
rect 1247 -17 1281 17
rect 1247 -85 1281 -51
rect 1405 51 1439 85
rect 1405 -17 1439 17
rect 1405 -85 1439 -51
rect 1563 51 1597 85
rect 1563 -17 1597 17
rect 1563 -85 1597 -51
rect 1721 51 1755 85
rect 1721 -17 1755 17
rect 1721 -85 1755 -51
rect 1879 51 1913 85
rect 1879 -17 1913 17
rect 1879 -85 1913 -51
rect 2037 51 2071 85
rect 2037 -17 2071 17
rect 2037 -85 2071 -51
rect 2195 51 2229 85
rect 2195 -17 2229 17
rect 2195 -85 2229 -51
rect 2353 51 2387 85
rect 2353 -17 2387 17
rect 2353 -85 2387 -51
rect 2511 51 2545 85
rect 2511 -17 2545 17
rect 2511 -85 2545 -51
rect 2669 51 2703 85
rect 2669 -17 2703 17
rect 2669 -85 2703 -51
rect 2827 51 2861 85
rect 2827 -17 2861 17
rect 2827 -85 2861 -51
rect 2985 51 3019 85
rect 2985 -17 3019 17
rect 2985 -85 3019 -51
rect 3143 51 3177 85
rect 3143 -17 3177 17
rect 3143 -85 3177 -51
rect -3177 -367 -3143 -333
rect -3177 -435 -3143 -401
rect -3177 -503 -3143 -469
rect -3019 -367 -2985 -333
rect -3019 -435 -2985 -401
rect -3019 -503 -2985 -469
rect -2861 -367 -2827 -333
rect -2861 -435 -2827 -401
rect -2861 -503 -2827 -469
rect -2703 -367 -2669 -333
rect -2703 -435 -2669 -401
rect -2703 -503 -2669 -469
rect -2545 -367 -2511 -333
rect -2545 -435 -2511 -401
rect -2545 -503 -2511 -469
rect -2387 -367 -2353 -333
rect -2387 -435 -2353 -401
rect -2387 -503 -2353 -469
rect -2229 -367 -2195 -333
rect -2229 -435 -2195 -401
rect -2229 -503 -2195 -469
rect -2071 -367 -2037 -333
rect -2071 -435 -2037 -401
rect -2071 -503 -2037 -469
rect -1913 -367 -1879 -333
rect -1913 -435 -1879 -401
rect -1913 -503 -1879 -469
rect -1755 -367 -1721 -333
rect -1755 -435 -1721 -401
rect -1755 -503 -1721 -469
rect -1597 -367 -1563 -333
rect -1597 -435 -1563 -401
rect -1597 -503 -1563 -469
rect -1439 -367 -1405 -333
rect -1439 -435 -1405 -401
rect -1439 -503 -1405 -469
rect -1281 -367 -1247 -333
rect -1281 -435 -1247 -401
rect -1281 -503 -1247 -469
rect -1123 -367 -1089 -333
rect -1123 -435 -1089 -401
rect -1123 -503 -1089 -469
rect -965 -367 -931 -333
rect -965 -435 -931 -401
rect -965 -503 -931 -469
rect -807 -367 -773 -333
rect -807 -435 -773 -401
rect -807 -503 -773 -469
rect -649 -367 -615 -333
rect -649 -435 -615 -401
rect -649 -503 -615 -469
rect -491 -367 -457 -333
rect -491 -435 -457 -401
rect -491 -503 -457 -469
rect -333 -367 -299 -333
rect -333 -435 -299 -401
rect -333 -503 -299 -469
rect -175 -367 -141 -333
rect -175 -435 -141 -401
rect -175 -503 -141 -469
rect -17 -367 17 -333
rect -17 -435 17 -401
rect -17 -503 17 -469
rect 141 -367 175 -333
rect 141 -435 175 -401
rect 141 -503 175 -469
rect 299 -367 333 -333
rect 299 -435 333 -401
rect 299 -503 333 -469
rect 457 -367 491 -333
rect 457 -435 491 -401
rect 457 -503 491 -469
rect 615 -367 649 -333
rect 615 -435 649 -401
rect 615 -503 649 -469
rect 773 -367 807 -333
rect 773 -435 807 -401
rect 773 -503 807 -469
rect 931 -367 965 -333
rect 931 -435 965 -401
rect 931 -503 965 -469
rect 1089 -367 1123 -333
rect 1089 -435 1123 -401
rect 1089 -503 1123 -469
rect 1247 -367 1281 -333
rect 1247 -435 1281 -401
rect 1247 -503 1281 -469
rect 1405 -367 1439 -333
rect 1405 -435 1439 -401
rect 1405 -503 1439 -469
rect 1563 -367 1597 -333
rect 1563 -435 1597 -401
rect 1563 -503 1597 -469
rect 1721 -367 1755 -333
rect 1721 -435 1755 -401
rect 1721 -503 1755 -469
rect 1879 -367 1913 -333
rect 1879 -435 1913 -401
rect 1879 -503 1913 -469
rect 2037 -367 2071 -333
rect 2037 -435 2071 -401
rect 2037 -503 2071 -469
rect 2195 -367 2229 -333
rect 2195 -435 2229 -401
rect 2195 -503 2229 -469
rect 2353 -367 2387 -333
rect 2353 -435 2387 -401
rect 2353 -503 2387 -469
rect 2511 -367 2545 -333
rect 2511 -435 2545 -401
rect 2511 -503 2545 -469
rect 2669 -367 2703 -333
rect 2669 -435 2703 -401
rect 2669 -503 2703 -469
rect 2827 -367 2861 -333
rect 2827 -435 2861 -401
rect 2827 -503 2861 -469
rect 2985 -367 3019 -333
rect 2985 -435 3019 -401
rect 2985 -503 3019 -469
rect 3143 -367 3177 -333
rect 3143 -435 3177 -401
rect 3143 -503 3177 -469
<< mvpsubdiff >>
rect -3323 728 3323 740
rect -3323 694 -3213 728
rect -3179 694 -3145 728
rect -3111 694 -3077 728
rect -3043 694 -3009 728
rect -2975 694 -2941 728
rect -2907 694 -2873 728
rect -2839 694 -2805 728
rect -2771 694 -2737 728
rect -2703 694 -2669 728
rect -2635 694 -2601 728
rect -2567 694 -2533 728
rect -2499 694 -2465 728
rect -2431 694 -2397 728
rect -2363 694 -2329 728
rect -2295 694 -2261 728
rect -2227 694 -2193 728
rect -2159 694 -2125 728
rect -2091 694 -2057 728
rect -2023 694 -1989 728
rect -1955 694 -1921 728
rect -1887 694 -1853 728
rect -1819 694 -1785 728
rect -1751 694 -1717 728
rect -1683 694 -1649 728
rect -1615 694 -1581 728
rect -1547 694 -1513 728
rect -1479 694 -1445 728
rect -1411 694 -1377 728
rect -1343 694 -1309 728
rect -1275 694 -1241 728
rect -1207 694 -1173 728
rect -1139 694 -1105 728
rect -1071 694 -1037 728
rect -1003 694 -969 728
rect -935 694 -901 728
rect -867 694 -833 728
rect -799 694 -765 728
rect -731 694 -697 728
rect -663 694 -629 728
rect -595 694 -561 728
rect -527 694 -493 728
rect -459 694 -425 728
rect -391 694 -357 728
rect -323 694 -289 728
rect -255 694 -221 728
rect -187 694 -153 728
rect -119 694 -85 728
rect -51 694 -17 728
rect 17 694 51 728
rect 85 694 119 728
rect 153 694 187 728
rect 221 694 255 728
rect 289 694 323 728
rect 357 694 391 728
rect 425 694 459 728
rect 493 694 527 728
rect 561 694 595 728
rect 629 694 663 728
rect 697 694 731 728
rect 765 694 799 728
rect 833 694 867 728
rect 901 694 935 728
rect 969 694 1003 728
rect 1037 694 1071 728
rect 1105 694 1139 728
rect 1173 694 1207 728
rect 1241 694 1275 728
rect 1309 694 1343 728
rect 1377 694 1411 728
rect 1445 694 1479 728
rect 1513 694 1547 728
rect 1581 694 1615 728
rect 1649 694 1683 728
rect 1717 694 1751 728
rect 1785 694 1819 728
rect 1853 694 1887 728
rect 1921 694 1955 728
rect 1989 694 2023 728
rect 2057 694 2091 728
rect 2125 694 2159 728
rect 2193 694 2227 728
rect 2261 694 2295 728
rect 2329 694 2363 728
rect 2397 694 2431 728
rect 2465 694 2499 728
rect 2533 694 2567 728
rect 2601 694 2635 728
rect 2669 694 2703 728
rect 2737 694 2771 728
rect 2805 694 2839 728
rect 2873 694 2907 728
rect 2941 694 2975 728
rect 3009 694 3043 728
rect 3077 694 3111 728
rect 3145 694 3179 728
rect 3213 694 3323 728
rect -3323 682 3323 694
rect -3323 629 -3265 682
rect -3323 595 -3311 629
rect -3277 595 -3265 629
rect 3265 629 3323 682
rect -3323 561 -3265 595
rect -3323 527 -3311 561
rect -3277 527 -3265 561
rect -3323 493 -3265 527
rect 3265 595 3277 629
rect 3311 595 3323 629
rect 3265 561 3323 595
rect 3265 527 3277 561
rect 3311 527 3323 561
rect -3323 459 -3311 493
rect -3277 459 -3265 493
rect -3323 425 -3265 459
rect -3323 391 -3311 425
rect -3277 391 -3265 425
rect -3323 357 -3265 391
rect -3323 323 -3311 357
rect -3277 323 -3265 357
rect -3323 289 -3265 323
rect 3265 493 3323 527
rect 3265 459 3277 493
rect 3311 459 3323 493
rect 3265 425 3323 459
rect 3265 391 3277 425
rect 3311 391 3323 425
rect 3265 357 3323 391
rect 3265 323 3277 357
rect 3311 323 3323 357
rect -3323 255 -3311 289
rect -3277 255 -3265 289
rect -3323 221 -3265 255
rect 3265 289 3323 323
rect 3265 255 3277 289
rect 3311 255 3323 289
rect -3323 187 -3311 221
rect -3277 187 -3265 221
rect 3265 221 3323 255
rect -3323 153 -3265 187
rect -3323 119 -3311 153
rect -3277 119 -3265 153
rect -3323 85 -3265 119
rect 3265 187 3277 221
rect 3311 187 3323 221
rect 3265 153 3323 187
rect 3265 119 3277 153
rect 3311 119 3323 153
rect -3323 51 -3311 85
rect -3277 51 -3265 85
rect -3323 17 -3265 51
rect -3323 -17 -3311 17
rect -3277 -17 -3265 17
rect -3323 -51 -3265 -17
rect -3323 -85 -3311 -51
rect -3277 -85 -3265 -51
rect -3323 -119 -3265 -85
rect 3265 85 3323 119
rect 3265 51 3277 85
rect 3311 51 3323 85
rect 3265 17 3323 51
rect 3265 -17 3277 17
rect 3311 -17 3323 17
rect 3265 -51 3323 -17
rect 3265 -85 3277 -51
rect 3311 -85 3323 -51
rect -3323 -153 -3311 -119
rect -3277 -153 -3265 -119
rect -3323 -187 -3265 -153
rect -3323 -221 -3311 -187
rect -3277 -221 -3265 -187
rect 3265 -119 3323 -85
rect 3265 -153 3277 -119
rect 3311 -153 3323 -119
rect 3265 -187 3323 -153
rect -3323 -255 -3265 -221
rect 3265 -221 3277 -187
rect 3311 -221 3323 -187
rect -3323 -289 -3311 -255
rect -3277 -289 -3265 -255
rect -3323 -323 -3265 -289
rect 3265 -255 3323 -221
rect 3265 -289 3277 -255
rect 3311 -289 3323 -255
rect -3323 -357 -3311 -323
rect -3277 -357 -3265 -323
rect -3323 -391 -3265 -357
rect -3323 -425 -3311 -391
rect -3277 -425 -3265 -391
rect -3323 -459 -3265 -425
rect -3323 -493 -3311 -459
rect -3277 -493 -3265 -459
rect -3323 -527 -3265 -493
rect 3265 -323 3323 -289
rect 3265 -357 3277 -323
rect 3311 -357 3323 -323
rect 3265 -391 3323 -357
rect 3265 -425 3277 -391
rect 3311 -425 3323 -391
rect 3265 -459 3323 -425
rect 3265 -493 3277 -459
rect 3311 -493 3323 -459
rect -3323 -561 -3311 -527
rect -3277 -561 -3265 -527
rect -3323 -595 -3265 -561
rect -3323 -629 -3311 -595
rect -3277 -629 -3265 -595
rect 3265 -527 3323 -493
rect 3265 -561 3277 -527
rect 3311 -561 3323 -527
rect 3265 -595 3323 -561
rect -3323 -682 -3265 -629
rect 3265 -629 3277 -595
rect 3311 -629 3323 -595
rect 3265 -682 3323 -629
rect -3323 -694 3323 -682
rect -3323 -728 -3213 -694
rect -3179 -728 -3145 -694
rect -3111 -728 -3077 -694
rect -3043 -728 -3009 -694
rect -2975 -728 -2941 -694
rect -2907 -728 -2873 -694
rect -2839 -728 -2805 -694
rect -2771 -728 -2737 -694
rect -2703 -728 -2669 -694
rect -2635 -728 -2601 -694
rect -2567 -728 -2533 -694
rect -2499 -728 -2465 -694
rect -2431 -728 -2397 -694
rect -2363 -728 -2329 -694
rect -2295 -728 -2261 -694
rect -2227 -728 -2193 -694
rect -2159 -728 -2125 -694
rect -2091 -728 -2057 -694
rect -2023 -728 -1989 -694
rect -1955 -728 -1921 -694
rect -1887 -728 -1853 -694
rect -1819 -728 -1785 -694
rect -1751 -728 -1717 -694
rect -1683 -728 -1649 -694
rect -1615 -728 -1581 -694
rect -1547 -728 -1513 -694
rect -1479 -728 -1445 -694
rect -1411 -728 -1377 -694
rect -1343 -728 -1309 -694
rect -1275 -728 -1241 -694
rect -1207 -728 -1173 -694
rect -1139 -728 -1105 -694
rect -1071 -728 -1037 -694
rect -1003 -728 -969 -694
rect -935 -728 -901 -694
rect -867 -728 -833 -694
rect -799 -728 -765 -694
rect -731 -728 -697 -694
rect -663 -728 -629 -694
rect -595 -728 -561 -694
rect -527 -728 -493 -694
rect -459 -728 -425 -694
rect -391 -728 -357 -694
rect -323 -728 -289 -694
rect -255 -728 -221 -694
rect -187 -728 -153 -694
rect -119 -728 -85 -694
rect -51 -728 -17 -694
rect 17 -728 51 -694
rect 85 -728 119 -694
rect 153 -728 187 -694
rect 221 -728 255 -694
rect 289 -728 323 -694
rect 357 -728 391 -694
rect 425 -728 459 -694
rect 493 -728 527 -694
rect 561 -728 595 -694
rect 629 -728 663 -694
rect 697 -728 731 -694
rect 765 -728 799 -694
rect 833 -728 867 -694
rect 901 -728 935 -694
rect 969 -728 1003 -694
rect 1037 -728 1071 -694
rect 1105 -728 1139 -694
rect 1173 -728 1207 -694
rect 1241 -728 1275 -694
rect 1309 -728 1343 -694
rect 1377 -728 1411 -694
rect 1445 -728 1479 -694
rect 1513 -728 1547 -694
rect 1581 -728 1615 -694
rect 1649 -728 1683 -694
rect 1717 -728 1751 -694
rect 1785 -728 1819 -694
rect 1853 -728 1887 -694
rect 1921 -728 1955 -694
rect 1989 -728 2023 -694
rect 2057 -728 2091 -694
rect 2125 -728 2159 -694
rect 2193 -728 2227 -694
rect 2261 -728 2295 -694
rect 2329 -728 2363 -694
rect 2397 -728 2431 -694
rect 2465 -728 2499 -694
rect 2533 -728 2567 -694
rect 2601 -728 2635 -694
rect 2669 -728 2703 -694
rect 2737 -728 2771 -694
rect 2805 -728 2839 -694
rect 2873 -728 2907 -694
rect 2941 -728 2975 -694
rect 3009 -728 3043 -694
rect 3077 -728 3111 -694
rect 3145 -728 3179 -694
rect 3213 -728 3323 -694
rect -3323 -740 3323 -728
<< mvpsubdiffcont >>
rect -3213 694 -3179 728
rect -3145 694 -3111 728
rect -3077 694 -3043 728
rect -3009 694 -2975 728
rect -2941 694 -2907 728
rect -2873 694 -2839 728
rect -2805 694 -2771 728
rect -2737 694 -2703 728
rect -2669 694 -2635 728
rect -2601 694 -2567 728
rect -2533 694 -2499 728
rect -2465 694 -2431 728
rect -2397 694 -2363 728
rect -2329 694 -2295 728
rect -2261 694 -2227 728
rect -2193 694 -2159 728
rect -2125 694 -2091 728
rect -2057 694 -2023 728
rect -1989 694 -1955 728
rect -1921 694 -1887 728
rect -1853 694 -1819 728
rect -1785 694 -1751 728
rect -1717 694 -1683 728
rect -1649 694 -1615 728
rect -1581 694 -1547 728
rect -1513 694 -1479 728
rect -1445 694 -1411 728
rect -1377 694 -1343 728
rect -1309 694 -1275 728
rect -1241 694 -1207 728
rect -1173 694 -1139 728
rect -1105 694 -1071 728
rect -1037 694 -1003 728
rect -969 694 -935 728
rect -901 694 -867 728
rect -833 694 -799 728
rect -765 694 -731 728
rect -697 694 -663 728
rect -629 694 -595 728
rect -561 694 -527 728
rect -493 694 -459 728
rect -425 694 -391 728
rect -357 694 -323 728
rect -289 694 -255 728
rect -221 694 -187 728
rect -153 694 -119 728
rect -85 694 -51 728
rect -17 694 17 728
rect 51 694 85 728
rect 119 694 153 728
rect 187 694 221 728
rect 255 694 289 728
rect 323 694 357 728
rect 391 694 425 728
rect 459 694 493 728
rect 527 694 561 728
rect 595 694 629 728
rect 663 694 697 728
rect 731 694 765 728
rect 799 694 833 728
rect 867 694 901 728
rect 935 694 969 728
rect 1003 694 1037 728
rect 1071 694 1105 728
rect 1139 694 1173 728
rect 1207 694 1241 728
rect 1275 694 1309 728
rect 1343 694 1377 728
rect 1411 694 1445 728
rect 1479 694 1513 728
rect 1547 694 1581 728
rect 1615 694 1649 728
rect 1683 694 1717 728
rect 1751 694 1785 728
rect 1819 694 1853 728
rect 1887 694 1921 728
rect 1955 694 1989 728
rect 2023 694 2057 728
rect 2091 694 2125 728
rect 2159 694 2193 728
rect 2227 694 2261 728
rect 2295 694 2329 728
rect 2363 694 2397 728
rect 2431 694 2465 728
rect 2499 694 2533 728
rect 2567 694 2601 728
rect 2635 694 2669 728
rect 2703 694 2737 728
rect 2771 694 2805 728
rect 2839 694 2873 728
rect 2907 694 2941 728
rect 2975 694 3009 728
rect 3043 694 3077 728
rect 3111 694 3145 728
rect 3179 694 3213 728
rect -3311 595 -3277 629
rect -3311 527 -3277 561
rect 3277 595 3311 629
rect 3277 527 3311 561
rect -3311 459 -3277 493
rect -3311 391 -3277 425
rect -3311 323 -3277 357
rect 3277 459 3311 493
rect 3277 391 3311 425
rect 3277 323 3311 357
rect -3311 255 -3277 289
rect 3277 255 3311 289
rect -3311 187 -3277 221
rect -3311 119 -3277 153
rect 3277 187 3311 221
rect 3277 119 3311 153
rect -3311 51 -3277 85
rect -3311 -17 -3277 17
rect -3311 -85 -3277 -51
rect 3277 51 3311 85
rect 3277 -17 3311 17
rect 3277 -85 3311 -51
rect -3311 -153 -3277 -119
rect -3311 -221 -3277 -187
rect 3277 -153 3311 -119
rect 3277 -221 3311 -187
rect -3311 -289 -3277 -255
rect 3277 -289 3311 -255
rect -3311 -357 -3277 -323
rect -3311 -425 -3277 -391
rect -3311 -493 -3277 -459
rect 3277 -357 3311 -323
rect 3277 -425 3311 -391
rect 3277 -493 3311 -459
rect -3311 -561 -3277 -527
rect -3311 -629 -3277 -595
rect 3277 -561 3311 -527
rect 3277 -629 3311 -595
rect -3213 -728 -3179 -694
rect -3145 -728 -3111 -694
rect -3077 -728 -3043 -694
rect -3009 -728 -2975 -694
rect -2941 -728 -2907 -694
rect -2873 -728 -2839 -694
rect -2805 -728 -2771 -694
rect -2737 -728 -2703 -694
rect -2669 -728 -2635 -694
rect -2601 -728 -2567 -694
rect -2533 -728 -2499 -694
rect -2465 -728 -2431 -694
rect -2397 -728 -2363 -694
rect -2329 -728 -2295 -694
rect -2261 -728 -2227 -694
rect -2193 -728 -2159 -694
rect -2125 -728 -2091 -694
rect -2057 -728 -2023 -694
rect -1989 -728 -1955 -694
rect -1921 -728 -1887 -694
rect -1853 -728 -1819 -694
rect -1785 -728 -1751 -694
rect -1717 -728 -1683 -694
rect -1649 -728 -1615 -694
rect -1581 -728 -1547 -694
rect -1513 -728 -1479 -694
rect -1445 -728 -1411 -694
rect -1377 -728 -1343 -694
rect -1309 -728 -1275 -694
rect -1241 -728 -1207 -694
rect -1173 -728 -1139 -694
rect -1105 -728 -1071 -694
rect -1037 -728 -1003 -694
rect -969 -728 -935 -694
rect -901 -728 -867 -694
rect -833 -728 -799 -694
rect -765 -728 -731 -694
rect -697 -728 -663 -694
rect -629 -728 -595 -694
rect -561 -728 -527 -694
rect -493 -728 -459 -694
rect -425 -728 -391 -694
rect -357 -728 -323 -694
rect -289 -728 -255 -694
rect -221 -728 -187 -694
rect -153 -728 -119 -694
rect -85 -728 -51 -694
rect -17 -728 17 -694
rect 51 -728 85 -694
rect 119 -728 153 -694
rect 187 -728 221 -694
rect 255 -728 289 -694
rect 323 -728 357 -694
rect 391 -728 425 -694
rect 459 -728 493 -694
rect 527 -728 561 -694
rect 595 -728 629 -694
rect 663 -728 697 -694
rect 731 -728 765 -694
rect 799 -728 833 -694
rect 867 -728 901 -694
rect 935 -728 969 -694
rect 1003 -728 1037 -694
rect 1071 -728 1105 -694
rect 1139 -728 1173 -694
rect 1207 -728 1241 -694
rect 1275 -728 1309 -694
rect 1343 -728 1377 -694
rect 1411 -728 1445 -694
rect 1479 -728 1513 -694
rect 1547 -728 1581 -694
rect 1615 -728 1649 -694
rect 1683 -728 1717 -694
rect 1751 -728 1785 -694
rect 1819 -728 1853 -694
rect 1887 -728 1921 -694
rect 1955 -728 1989 -694
rect 2023 -728 2057 -694
rect 2091 -728 2125 -694
rect 2159 -728 2193 -694
rect 2227 -728 2261 -694
rect 2295 -728 2329 -694
rect 2363 -728 2397 -694
rect 2431 -728 2465 -694
rect 2499 -728 2533 -694
rect 2567 -728 2601 -694
rect 2635 -728 2669 -694
rect 2703 -728 2737 -694
rect 2771 -728 2805 -694
rect 2839 -728 2873 -694
rect 2907 -728 2941 -694
rect 2975 -728 3009 -694
rect 3043 -728 3077 -694
rect 3111 -728 3145 -694
rect 3179 -728 3213 -694
<< poly >>
rect -3131 590 -3031 606
rect -3131 556 -3098 590
rect -3064 556 -3031 590
rect -3131 518 -3031 556
rect -2973 590 -2873 606
rect -2973 556 -2940 590
rect -2906 556 -2873 590
rect -2973 518 -2873 556
rect -2815 590 -2715 606
rect -2815 556 -2782 590
rect -2748 556 -2715 590
rect -2815 518 -2715 556
rect -2657 590 -2557 606
rect -2657 556 -2624 590
rect -2590 556 -2557 590
rect -2657 518 -2557 556
rect -2499 590 -2399 606
rect -2499 556 -2466 590
rect -2432 556 -2399 590
rect -2499 518 -2399 556
rect -2341 590 -2241 606
rect -2341 556 -2308 590
rect -2274 556 -2241 590
rect -2341 518 -2241 556
rect -2183 590 -2083 606
rect -2183 556 -2150 590
rect -2116 556 -2083 590
rect -2183 518 -2083 556
rect -2025 590 -1925 606
rect -2025 556 -1992 590
rect -1958 556 -1925 590
rect -2025 518 -1925 556
rect -1867 590 -1767 606
rect -1867 556 -1834 590
rect -1800 556 -1767 590
rect -1867 518 -1767 556
rect -1709 590 -1609 606
rect -1709 556 -1676 590
rect -1642 556 -1609 590
rect -1709 518 -1609 556
rect -1551 590 -1451 606
rect -1551 556 -1518 590
rect -1484 556 -1451 590
rect -1551 518 -1451 556
rect -1393 590 -1293 606
rect -1393 556 -1360 590
rect -1326 556 -1293 590
rect -1393 518 -1293 556
rect -1235 590 -1135 606
rect -1235 556 -1202 590
rect -1168 556 -1135 590
rect -1235 518 -1135 556
rect -1077 590 -977 606
rect -1077 556 -1044 590
rect -1010 556 -977 590
rect -1077 518 -977 556
rect -919 590 -819 606
rect -919 556 -886 590
rect -852 556 -819 590
rect -919 518 -819 556
rect -761 590 -661 606
rect -761 556 -728 590
rect -694 556 -661 590
rect -761 518 -661 556
rect -603 590 -503 606
rect -603 556 -570 590
rect -536 556 -503 590
rect -603 518 -503 556
rect -445 590 -345 606
rect -445 556 -412 590
rect -378 556 -345 590
rect -445 518 -345 556
rect -287 590 -187 606
rect -287 556 -254 590
rect -220 556 -187 590
rect -287 518 -187 556
rect -129 590 -29 606
rect -129 556 -96 590
rect -62 556 -29 590
rect -129 518 -29 556
rect 29 590 129 606
rect 29 556 62 590
rect 96 556 129 590
rect 29 518 129 556
rect 187 590 287 606
rect 187 556 220 590
rect 254 556 287 590
rect 187 518 287 556
rect 345 590 445 606
rect 345 556 378 590
rect 412 556 445 590
rect 345 518 445 556
rect 503 590 603 606
rect 503 556 536 590
rect 570 556 603 590
rect 503 518 603 556
rect 661 590 761 606
rect 661 556 694 590
rect 728 556 761 590
rect 661 518 761 556
rect 819 590 919 606
rect 819 556 852 590
rect 886 556 919 590
rect 819 518 919 556
rect 977 590 1077 606
rect 977 556 1010 590
rect 1044 556 1077 590
rect 977 518 1077 556
rect 1135 590 1235 606
rect 1135 556 1168 590
rect 1202 556 1235 590
rect 1135 518 1235 556
rect 1293 590 1393 606
rect 1293 556 1326 590
rect 1360 556 1393 590
rect 1293 518 1393 556
rect 1451 590 1551 606
rect 1451 556 1484 590
rect 1518 556 1551 590
rect 1451 518 1551 556
rect 1609 590 1709 606
rect 1609 556 1642 590
rect 1676 556 1709 590
rect 1609 518 1709 556
rect 1767 590 1867 606
rect 1767 556 1800 590
rect 1834 556 1867 590
rect 1767 518 1867 556
rect 1925 590 2025 606
rect 1925 556 1958 590
rect 1992 556 2025 590
rect 1925 518 2025 556
rect 2083 590 2183 606
rect 2083 556 2116 590
rect 2150 556 2183 590
rect 2083 518 2183 556
rect 2241 590 2341 606
rect 2241 556 2274 590
rect 2308 556 2341 590
rect 2241 518 2341 556
rect 2399 590 2499 606
rect 2399 556 2432 590
rect 2466 556 2499 590
rect 2399 518 2499 556
rect 2557 590 2657 606
rect 2557 556 2590 590
rect 2624 556 2657 590
rect 2557 518 2657 556
rect 2715 590 2815 606
rect 2715 556 2748 590
rect 2782 556 2815 590
rect 2715 518 2815 556
rect 2873 590 2973 606
rect 2873 556 2906 590
rect 2940 556 2973 590
rect 2873 518 2973 556
rect 3031 590 3131 606
rect 3031 556 3064 590
rect 3098 556 3131 590
rect 3031 518 3131 556
rect -3131 280 -3031 318
rect -3131 246 -3098 280
rect -3064 246 -3031 280
rect -3131 230 -3031 246
rect -2973 280 -2873 318
rect -2973 246 -2940 280
rect -2906 246 -2873 280
rect -2973 230 -2873 246
rect -2815 280 -2715 318
rect -2815 246 -2782 280
rect -2748 246 -2715 280
rect -2815 230 -2715 246
rect -2657 280 -2557 318
rect -2657 246 -2624 280
rect -2590 246 -2557 280
rect -2657 230 -2557 246
rect -2499 280 -2399 318
rect -2499 246 -2466 280
rect -2432 246 -2399 280
rect -2499 230 -2399 246
rect -2341 280 -2241 318
rect -2341 246 -2308 280
rect -2274 246 -2241 280
rect -2341 230 -2241 246
rect -2183 280 -2083 318
rect -2183 246 -2150 280
rect -2116 246 -2083 280
rect -2183 230 -2083 246
rect -2025 280 -1925 318
rect -2025 246 -1992 280
rect -1958 246 -1925 280
rect -2025 230 -1925 246
rect -1867 280 -1767 318
rect -1867 246 -1834 280
rect -1800 246 -1767 280
rect -1867 230 -1767 246
rect -1709 280 -1609 318
rect -1709 246 -1676 280
rect -1642 246 -1609 280
rect -1709 230 -1609 246
rect -1551 280 -1451 318
rect -1551 246 -1518 280
rect -1484 246 -1451 280
rect -1551 230 -1451 246
rect -1393 280 -1293 318
rect -1393 246 -1360 280
rect -1326 246 -1293 280
rect -1393 230 -1293 246
rect -1235 280 -1135 318
rect -1235 246 -1202 280
rect -1168 246 -1135 280
rect -1235 230 -1135 246
rect -1077 280 -977 318
rect -1077 246 -1044 280
rect -1010 246 -977 280
rect -1077 230 -977 246
rect -919 280 -819 318
rect -919 246 -886 280
rect -852 246 -819 280
rect -919 230 -819 246
rect -761 280 -661 318
rect -761 246 -728 280
rect -694 246 -661 280
rect -761 230 -661 246
rect -603 280 -503 318
rect -603 246 -570 280
rect -536 246 -503 280
rect -603 230 -503 246
rect -445 280 -345 318
rect -445 246 -412 280
rect -378 246 -345 280
rect -445 230 -345 246
rect -287 280 -187 318
rect -287 246 -254 280
rect -220 246 -187 280
rect -287 230 -187 246
rect -129 280 -29 318
rect -129 246 -96 280
rect -62 246 -29 280
rect -129 230 -29 246
rect 29 280 129 318
rect 29 246 62 280
rect 96 246 129 280
rect 29 230 129 246
rect 187 280 287 318
rect 187 246 220 280
rect 254 246 287 280
rect 187 230 287 246
rect 345 280 445 318
rect 345 246 378 280
rect 412 246 445 280
rect 345 230 445 246
rect 503 280 603 318
rect 503 246 536 280
rect 570 246 603 280
rect 503 230 603 246
rect 661 280 761 318
rect 661 246 694 280
rect 728 246 761 280
rect 661 230 761 246
rect 819 280 919 318
rect 819 246 852 280
rect 886 246 919 280
rect 819 230 919 246
rect 977 280 1077 318
rect 977 246 1010 280
rect 1044 246 1077 280
rect 977 230 1077 246
rect 1135 280 1235 318
rect 1135 246 1168 280
rect 1202 246 1235 280
rect 1135 230 1235 246
rect 1293 280 1393 318
rect 1293 246 1326 280
rect 1360 246 1393 280
rect 1293 230 1393 246
rect 1451 280 1551 318
rect 1451 246 1484 280
rect 1518 246 1551 280
rect 1451 230 1551 246
rect 1609 280 1709 318
rect 1609 246 1642 280
rect 1676 246 1709 280
rect 1609 230 1709 246
rect 1767 280 1867 318
rect 1767 246 1800 280
rect 1834 246 1867 280
rect 1767 230 1867 246
rect 1925 280 2025 318
rect 1925 246 1958 280
rect 1992 246 2025 280
rect 1925 230 2025 246
rect 2083 280 2183 318
rect 2083 246 2116 280
rect 2150 246 2183 280
rect 2083 230 2183 246
rect 2241 280 2341 318
rect 2241 246 2274 280
rect 2308 246 2341 280
rect 2241 230 2341 246
rect 2399 280 2499 318
rect 2399 246 2432 280
rect 2466 246 2499 280
rect 2399 230 2499 246
rect 2557 280 2657 318
rect 2557 246 2590 280
rect 2624 246 2657 280
rect 2557 230 2657 246
rect 2715 280 2815 318
rect 2715 246 2748 280
rect 2782 246 2815 280
rect 2715 230 2815 246
rect 2873 280 2973 318
rect 2873 246 2906 280
rect 2940 246 2973 280
rect 2873 230 2973 246
rect 3031 280 3131 318
rect 3031 246 3064 280
rect 3098 246 3131 280
rect 3031 230 3131 246
rect -3131 172 -3031 188
rect -3131 138 -3098 172
rect -3064 138 -3031 172
rect -3131 100 -3031 138
rect -2973 172 -2873 188
rect -2973 138 -2940 172
rect -2906 138 -2873 172
rect -2973 100 -2873 138
rect -2815 172 -2715 188
rect -2815 138 -2782 172
rect -2748 138 -2715 172
rect -2815 100 -2715 138
rect -2657 172 -2557 188
rect -2657 138 -2624 172
rect -2590 138 -2557 172
rect -2657 100 -2557 138
rect -2499 172 -2399 188
rect -2499 138 -2466 172
rect -2432 138 -2399 172
rect -2499 100 -2399 138
rect -2341 172 -2241 188
rect -2341 138 -2308 172
rect -2274 138 -2241 172
rect -2341 100 -2241 138
rect -2183 172 -2083 188
rect -2183 138 -2150 172
rect -2116 138 -2083 172
rect -2183 100 -2083 138
rect -2025 172 -1925 188
rect -2025 138 -1992 172
rect -1958 138 -1925 172
rect -2025 100 -1925 138
rect -1867 172 -1767 188
rect -1867 138 -1834 172
rect -1800 138 -1767 172
rect -1867 100 -1767 138
rect -1709 172 -1609 188
rect -1709 138 -1676 172
rect -1642 138 -1609 172
rect -1709 100 -1609 138
rect -1551 172 -1451 188
rect -1551 138 -1518 172
rect -1484 138 -1451 172
rect -1551 100 -1451 138
rect -1393 172 -1293 188
rect -1393 138 -1360 172
rect -1326 138 -1293 172
rect -1393 100 -1293 138
rect -1235 172 -1135 188
rect -1235 138 -1202 172
rect -1168 138 -1135 172
rect -1235 100 -1135 138
rect -1077 172 -977 188
rect -1077 138 -1044 172
rect -1010 138 -977 172
rect -1077 100 -977 138
rect -919 172 -819 188
rect -919 138 -886 172
rect -852 138 -819 172
rect -919 100 -819 138
rect -761 172 -661 188
rect -761 138 -728 172
rect -694 138 -661 172
rect -761 100 -661 138
rect -603 172 -503 188
rect -603 138 -570 172
rect -536 138 -503 172
rect -603 100 -503 138
rect -445 172 -345 188
rect -445 138 -412 172
rect -378 138 -345 172
rect -445 100 -345 138
rect -287 172 -187 188
rect -287 138 -254 172
rect -220 138 -187 172
rect -287 100 -187 138
rect -129 172 -29 188
rect -129 138 -96 172
rect -62 138 -29 172
rect -129 100 -29 138
rect 29 172 129 188
rect 29 138 62 172
rect 96 138 129 172
rect 29 100 129 138
rect 187 172 287 188
rect 187 138 220 172
rect 254 138 287 172
rect 187 100 287 138
rect 345 172 445 188
rect 345 138 378 172
rect 412 138 445 172
rect 345 100 445 138
rect 503 172 603 188
rect 503 138 536 172
rect 570 138 603 172
rect 503 100 603 138
rect 661 172 761 188
rect 661 138 694 172
rect 728 138 761 172
rect 661 100 761 138
rect 819 172 919 188
rect 819 138 852 172
rect 886 138 919 172
rect 819 100 919 138
rect 977 172 1077 188
rect 977 138 1010 172
rect 1044 138 1077 172
rect 977 100 1077 138
rect 1135 172 1235 188
rect 1135 138 1168 172
rect 1202 138 1235 172
rect 1135 100 1235 138
rect 1293 172 1393 188
rect 1293 138 1326 172
rect 1360 138 1393 172
rect 1293 100 1393 138
rect 1451 172 1551 188
rect 1451 138 1484 172
rect 1518 138 1551 172
rect 1451 100 1551 138
rect 1609 172 1709 188
rect 1609 138 1642 172
rect 1676 138 1709 172
rect 1609 100 1709 138
rect 1767 172 1867 188
rect 1767 138 1800 172
rect 1834 138 1867 172
rect 1767 100 1867 138
rect 1925 172 2025 188
rect 1925 138 1958 172
rect 1992 138 2025 172
rect 1925 100 2025 138
rect 2083 172 2183 188
rect 2083 138 2116 172
rect 2150 138 2183 172
rect 2083 100 2183 138
rect 2241 172 2341 188
rect 2241 138 2274 172
rect 2308 138 2341 172
rect 2241 100 2341 138
rect 2399 172 2499 188
rect 2399 138 2432 172
rect 2466 138 2499 172
rect 2399 100 2499 138
rect 2557 172 2657 188
rect 2557 138 2590 172
rect 2624 138 2657 172
rect 2557 100 2657 138
rect 2715 172 2815 188
rect 2715 138 2748 172
rect 2782 138 2815 172
rect 2715 100 2815 138
rect 2873 172 2973 188
rect 2873 138 2906 172
rect 2940 138 2973 172
rect 2873 100 2973 138
rect 3031 172 3131 188
rect 3031 138 3064 172
rect 3098 138 3131 172
rect 3031 100 3131 138
rect -3131 -138 -3031 -100
rect -3131 -172 -3098 -138
rect -3064 -172 -3031 -138
rect -3131 -188 -3031 -172
rect -2973 -138 -2873 -100
rect -2973 -172 -2940 -138
rect -2906 -172 -2873 -138
rect -2973 -188 -2873 -172
rect -2815 -138 -2715 -100
rect -2815 -172 -2782 -138
rect -2748 -172 -2715 -138
rect -2815 -188 -2715 -172
rect -2657 -138 -2557 -100
rect -2657 -172 -2624 -138
rect -2590 -172 -2557 -138
rect -2657 -188 -2557 -172
rect -2499 -138 -2399 -100
rect -2499 -172 -2466 -138
rect -2432 -172 -2399 -138
rect -2499 -188 -2399 -172
rect -2341 -138 -2241 -100
rect -2341 -172 -2308 -138
rect -2274 -172 -2241 -138
rect -2341 -188 -2241 -172
rect -2183 -138 -2083 -100
rect -2183 -172 -2150 -138
rect -2116 -172 -2083 -138
rect -2183 -188 -2083 -172
rect -2025 -138 -1925 -100
rect -2025 -172 -1992 -138
rect -1958 -172 -1925 -138
rect -2025 -188 -1925 -172
rect -1867 -138 -1767 -100
rect -1867 -172 -1834 -138
rect -1800 -172 -1767 -138
rect -1867 -188 -1767 -172
rect -1709 -138 -1609 -100
rect -1709 -172 -1676 -138
rect -1642 -172 -1609 -138
rect -1709 -188 -1609 -172
rect -1551 -138 -1451 -100
rect -1551 -172 -1518 -138
rect -1484 -172 -1451 -138
rect -1551 -188 -1451 -172
rect -1393 -138 -1293 -100
rect -1393 -172 -1360 -138
rect -1326 -172 -1293 -138
rect -1393 -188 -1293 -172
rect -1235 -138 -1135 -100
rect -1235 -172 -1202 -138
rect -1168 -172 -1135 -138
rect -1235 -188 -1135 -172
rect -1077 -138 -977 -100
rect -1077 -172 -1044 -138
rect -1010 -172 -977 -138
rect -1077 -188 -977 -172
rect -919 -138 -819 -100
rect -919 -172 -886 -138
rect -852 -172 -819 -138
rect -919 -188 -819 -172
rect -761 -138 -661 -100
rect -761 -172 -728 -138
rect -694 -172 -661 -138
rect -761 -188 -661 -172
rect -603 -138 -503 -100
rect -603 -172 -570 -138
rect -536 -172 -503 -138
rect -603 -188 -503 -172
rect -445 -138 -345 -100
rect -445 -172 -412 -138
rect -378 -172 -345 -138
rect -445 -188 -345 -172
rect -287 -138 -187 -100
rect -287 -172 -254 -138
rect -220 -172 -187 -138
rect -287 -188 -187 -172
rect -129 -138 -29 -100
rect -129 -172 -96 -138
rect -62 -172 -29 -138
rect -129 -188 -29 -172
rect 29 -138 129 -100
rect 29 -172 62 -138
rect 96 -172 129 -138
rect 29 -188 129 -172
rect 187 -138 287 -100
rect 187 -172 220 -138
rect 254 -172 287 -138
rect 187 -188 287 -172
rect 345 -138 445 -100
rect 345 -172 378 -138
rect 412 -172 445 -138
rect 345 -188 445 -172
rect 503 -138 603 -100
rect 503 -172 536 -138
rect 570 -172 603 -138
rect 503 -188 603 -172
rect 661 -138 761 -100
rect 661 -172 694 -138
rect 728 -172 761 -138
rect 661 -188 761 -172
rect 819 -138 919 -100
rect 819 -172 852 -138
rect 886 -172 919 -138
rect 819 -188 919 -172
rect 977 -138 1077 -100
rect 977 -172 1010 -138
rect 1044 -172 1077 -138
rect 977 -188 1077 -172
rect 1135 -138 1235 -100
rect 1135 -172 1168 -138
rect 1202 -172 1235 -138
rect 1135 -188 1235 -172
rect 1293 -138 1393 -100
rect 1293 -172 1326 -138
rect 1360 -172 1393 -138
rect 1293 -188 1393 -172
rect 1451 -138 1551 -100
rect 1451 -172 1484 -138
rect 1518 -172 1551 -138
rect 1451 -188 1551 -172
rect 1609 -138 1709 -100
rect 1609 -172 1642 -138
rect 1676 -172 1709 -138
rect 1609 -188 1709 -172
rect 1767 -138 1867 -100
rect 1767 -172 1800 -138
rect 1834 -172 1867 -138
rect 1767 -188 1867 -172
rect 1925 -138 2025 -100
rect 1925 -172 1958 -138
rect 1992 -172 2025 -138
rect 1925 -188 2025 -172
rect 2083 -138 2183 -100
rect 2083 -172 2116 -138
rect 2150 -172 2183 -138
rect 2083 -188 2183 -172
rect 2241 -138 2341 -100
rect 2241 -172 2274 -138
rect 2308 -172 2341 -138
rect 2241 -188 2341 -172
rect 2399 -138 2499 -100
rect 2399 -172 2432 -138
rect 2466 -172 2499 -138
rect 2399 -188 2499 -172
rect 2557 -138 2657 -100
rect 2557 -172 2590 -138
rect 2624 -172 2657 -138
rect 2557 -188 2657 -172
rect 2715 -138 2815 -100
rect 2715 -172 2748 -138
rect 2782 -172 2815 -138
rect 2715 -188 2815 -172
rect 2873 -138 2973 -100
rect 2873 -172 2906 -138
rect 2940 -172 2973 -138
rect 2873 -188 2973 -172
rect 3031 -138 3131 -100
rect 3031 -172 3064 -138
rect 3098 -172 3131 -138
rect 3031 -188 3131 -172
rect -3131 -246 -3031 -230
rect -3131 -280 -3098 -246
rect -3064 -280 -3031 -246
rect -3131 -318 -3031 -280
rect -2973 -246 -2873 -230
rect -2973 -280 -2940 -246
rect -2906 -280 -2873 -246
rect -2973 -318 -2873 -280
rect -2815 -246 -2715 -230
rect -2815 -280 -2782 -246
rect -2748 -280 -2715 -246
rect -2815 -318 -2715 -280
rect -2657 -246 -2557 -230
rect -2657 -280 -2624 -246
rect -2590 -280 -2557 -246
rect -2657 -318 -2557 -280
rect -2499 -246 -2399 -230
rect -2499 -280 -2466 -246
rect -2432 -280 -2399 -246
rect -2499 -318 -2399 -280
rect -2341 -246 -2241 -230
rect -2341 -280 -2308 -246
rect -2274 -280 -2241 -246
rect -2341 -318 -2241 -280
rect -2183 -246 -2083 -230
rect -2183 -280 -2150 -246
rect -2116 -280 -2083 -246
rect -2183 -318 -2083 -280
rect -2025 -246 -1925 -230
rect -2025 -280 -1992 -246
rect -1958 -280 -1925 -246
rect -2025 -318 -1925 -280
rect -1867 -246 -1767 -230
rect -1867 -280 -1834 -246
rect -1800 -280 -1767 -246
rect -1867 -318 -1767 -280
rect -1709 -246 -1609 -230
rect -1709 -280 -1676 -246
rect -1642 -280 -1609 -246
rect -1709 -318 -1609 -280
rect -1551 -246 -1451 -230
rect -1551 -280 -1518 -246
rect -1484 -280 -1451 -246
rect -1551 -318 -1451 -280
rect -1393 -246 -1293 -230
rect -1393 -280 -1360 -246
rect -1326 -280 -1293 -246
rect -1393 -318 -1293 -280
rect -1235 -246 -1135 -230
rect -1235 -280 -1202 -246
rect -1168 -280 -1135 -246
rect -1235 -318 -1135 -280
rect -1077 -246 -977 -230
rect -1077 -280 -1044 -246
rect -1010 -280 -977 -246
rect -1077 -318 -977 -280
rect -919 -246 -819 -230
rect -919 -280 -886 -246
rect -852 -280 -819 -246
rect -919 -318 -819 -280
rect -761 -246 -661 -230
rect -761 -280 -728 -246
rect -694 -280 -661 -246
rect -761 -318 -661 -280
rect -603 -246 -503 -230
rect -603 -280 -570 -246
rect -536 -280 -503 -246
rect -603 -318 -503 -280
rect -445 -246 -345 -230
rect -445 -280 -412 -246
rect -378 -280 -345 -246
rect -445 -318 -345 -280
rect -287 -246 -187 -230
rect -287 -280 -254 -246
rect -220 -280 -187 -246
rect -287 -318 -187 -280
rect -129 -246 -29 -230
rect -129 -280 -96 -246
rect -62 -280 -29 -246
rect -129 -318 -29 -280
rect 29 -246 129 -230
rect 29 -280 62 -246
rect 96 -280 129 -246
rect 29 -318 129 -280
rect 187 -246 287 -230
rect 187 -280 220 -246
rect 254 -280 287 -246
rect 187 -318 287 -280
rect 345 -246 445 -230
rect 345 -280 378 -246
rect 412 -280 445 -246
rect 345 -318 445 -280
rect 503 -246 603 -230
rect 503 -280 536 -246
rect 570 -280 603 -246
rect 503 -318 603 -280
rect 661 -246 761 -230
rect 661 -280 694 -246
rect 728 -280 761 -246
rect 661 -318 761 -280
rect 819 -246 919 -230
rect 819 -280 852 -246
rect 886 -280 919 -246
rect 819 -318 919 -280
rect 977 -246 1077 -230
rect 977 -280 1010 -246
rect 1044 -280 1077 -246
rect 977 -318 1077 -280
rect 1135 -246 1235 -230
rect 1135 -280 1168 -246
rect 1202 -280 1235 -246
rect 1135 -318 1235 -280
rect 1293 -246 1393 -230
rect 1293 -280 1326 -246
rect 1360 -280 1393 -246
rect 1293 -318 1393 -280
rect 1451 -246 1551 -230
rect 1451 -280 1484 -246
rect 1518 -280 1551 -246
rect 1451 -318 1551 -280
rect 1609 -246 1709 -230
rect 1609 -280 1642 -246
rect 1676 -280 1709 -246
rect 1609 -318 1709 -280
rect 1767 -246 1867 -230
rect 1767 -280 1800 -246
rect 1834 -280 1867 -246
rect 1767 -318 1867 -280
rect 1925 -246 2025 -230
rect 1925 -280 1958 -246
rect 1992 -280 2025 -246
rect 1925 -318 2025 -280
rect 2083 -246 2183 -230
rect 2083 -280 2116 -246
rect 2150 -280 2183 -246
rect 2083 -318 2183 -280
rect 2241 -246 2341 -230
rect 2241 -280 2274 -246
rect 2308 -280 2341 -246
rect 2241 -318 2341 -280
rect 2399 -246 2499 -230
rect 2399 -280 2432 -246
rect 2466 -280 2499 -246
rect 2399 -318 2499 -280
rect 2557 -246 2657 -230
rect 2557 -280 2590 -246
rect 2624 -280 2657 -246
rect 2557 -318 2657 -280
rect 2715 -246 2815 -230
rect 2715 -280 2748 -246
rect 2782 -280 2815 -246
rect 2715 -318 2815 -280
rect 2873 -246 2973 -230
rect 2873 -280 2906 -246
rect 2940 -280 2973 -246
rect 2873 -318 2973 -280
rect 3031 -246 3131 -230
rect 3031 -280 3064 -246
rect 3098 -280 3131 -246
rect 3031 -318 3131 -280
rect -3131 -556 -3031 -518
rect -3131 -590 -3098 -556
rect -3064 -590 -3031 -556
rect -3131 -606 -3031 -590
rect -2973 -556 -2873 -518
rect -2973 -590 -2940 -556
rect -2906 -590 -2873 -556
rect -2973 -606 -2873 -590
rect -2815 -556 -2715 -518
rect -2815 -590 -2782 -556
rect -2748 -590 -2715 -556
rect -2815 -606 -2715 -590
rect -2657 -556 -2557 -518
rect -2657 -590 -2624 -556
rect -2590 -590 -2557 -556
rect -2657 -606 -2557 -590
rect -2499 -556 -2399 -518
rect -2499 -590 -2466 -556
rect -2432 -590 -2399 -556
rect -2499 -606 -2399 -590
rect -2341 -556 -2241 -518
rect -2341 -590 -2308 -556
rect -2274 -590 -2241 -556
rect -2341 -606 -2241 -590
rect -2183 -556 -2083 -518
rect -2183 -590 -2150 -556
rect -2116 -590 -2083 -556
rect -2183 -606 -2083 -590
rect -2025 -556 -1925 -518
rect -2025 -590 -1992 -556
rect -1958 -590 -1925 -556
rect -2025 -606 -1925 -590
rect -1867 -556 -1767 -518
rect -1867 -590 -1834 -556
rect -1800 -590 -1767 -556
rect -1867 -606 -1767 -590
rect -1709 -556 -1609 -518
rect -1709 -590 -1676 -556
rect -1642 -590 -1609 -556
rect -1709 -606 -1609 -590
rect -1551 -556 -1451 -518
rect -1551 -590 -1518 -556
rect -1484 -590 -1451 -556
rect -1551 -606 -1451 -590
rect -1393 -556 -1293 -518
rect -1393 -590 -1360 -556
rect -1326 -590 -1293 -556
rect -1393 -606 -1293 -590
rect -1235 -556 -1135 -518
rect -1235 -590 -1202 -556
rect -1168 -590 -1135 -556
rect -1235 -606 -1135 -590
rect -1077 -556 -977 -518
rect -1077 -590 -1044 -556
rect -1010 -590 -977 -556
rect -1077 -606 -977 -590
rect -919 -556 -819 -518
rect -919 -590 -886 -556
rect -852 -590 -819 -556
rect -919 -606 -819 -590
rect -761 -556 -661 -518
rect -761 -590 -728 -556
rect -694 -590 -661 -556
rect -761 -606 -661 -590
rect -603 -556 -503 -518
rect -603 -590 -570 -556
rect -536 -590 -503 -556
rect -603 -606 -503 -590
rect -445 -556 -345 -518
rect -445 -590 -412 -556
rect -378 -590 -345 -556
rect -445 -606 -345 -590
rect -287 -556 -187 -518
rect -287 -590 -254 -556
rect -220 -590 -187 -556
rect -287 -606 -187 -590
rect -129 -556 -29 -518
rect -129 -590 -96 -556
rect -62 -590 -29 -556
rect -129 -606 -29 -590
rect 29 -556 129 -518
rect 29 -590 62 -556
rect 96 -590 129 -556
rect 29 -606 129 -590
rect 187 -556 287 -518
rect 187 -590 220 -556
rect 254 -590 287 -556
rect 187 -606 287 -590
rect 345 -556 445 -518
rect 345 -590 378 -556
rect 412 -590 445 -556
rect 345 -606 445 -590
rect 503 -556 603 -518
rect 503 -590 536 -556
rect 570 -590 603 -556
rect 503 -606 603 -590
rect 661 -556 761 -518
rect 661 -590 694 -556
rect 728 -590 761 -556
rect 661 -606 761 -590
rect 819 -556 919 -518
rect 819 -590 852 -556
rect 886 -590 919 -556
rect 819 -606 919 -590
rect 977 -556 1077 -518
rect 977 -590 1010 -556
rect 1044 -590 1077 -556
rect 977 -606 1077 -590
rect 1135 -556 1235 -518
rect 1135 -590 1168 -556
rect 1202 -590 1235 -556
rect 1135 -606 1235 -590
rect 1293 -556 1393 -518
rect 1293 -590 1326 -556
rect 1360 -590 1393 -556
rect 1293 -606 1393 -590
rect 1451 -556 1551 -518
rect 1451 -590 1484 -556
rect 1518 -590 1551 -556
rect 1451 -606 1551 -590
rect 1609 -556 1709 -518
rect 1609 -590 1642 -556
rect 1676 -590 1709 -556
rect 1609 -606 1709 -590
rect 1767 -556 1867 -518
rect 1767 -590 1800 -556
rect 1834 -590 1867 -556
rect 1767 -606 1867 -590
rect 1925 -556 2025 -518
rect 1925 -590 1958 -556
rect 1992 -590 2025 -556
rect 1925 -606 2025 -590
rect 2083 -556 2183 -518
rect 2083 -590 2116 -556
rect 2150 -590 2183 -556
rect 2083 -606 2183 -590
rect 2241 -556 2341 -518
rect 2241 -590 2274 -556
rect 2308 -590 2341 -556
rect 2241 -606 2341 -590
rect 2399 -556 2499 -518
rect 2399 -590 2432 -556
rect 2466 -590 2499 -556
rect 2399 -606 2499 -590
rect 2557 -556 2657 -518
rect 2557 -590 2590 -556
rect 2624 -590 2657 -556
rect 2557 -606 2657 -590
rect 2715 -556 2815 -518
rect 2715 -590 2748 -556
rect 2782 -590 2815 -556
rect 2715 -606 2815 -590
rect 2873 -556 2973 -518
rect 2873 -590 2906 -556
rect 2940 -590 2973 -556
rect 2873 -606 2973 -590
rect 3031 -556 3131 -518
rect 3031 -590 3064 -556
rect 3098 -590 3131 -556
rect 3031 -606 3131 -590
<< polycont >>
rect -3098 556 -3064 590
rect -2940 556 -2906 590
rect -2782 556 -2748 590
rect -2624 556 -2590 590
rect -2466 556 -2432 590
rect -2308 556 -2274 590
rect -2150 556 -2116 590
rect -1992 556 -1958 590
rect -1834 556 -1800 590
rect -1676 556 -1642 590
rect -1518 556 -1484 590
rect -1360 556 -1326 590
rect -1202 556 -1168 590
rect -1044 556 -1010 590
rect -886 556 -852 590
rect -728 556 -694 590
rect -570 556 -536 590
rect -412 556 -378 590
rect -254 556 -220 590
rect -96 556 -62 590
rect 62 556 96 590
rect 220 556 254 590
rect 378 556 412 590
rect 536 556 570 590
rect 694 556 728 590
rect 852 556 886 590
rect 1010 556 1044 590
rect 1168 556 1202 590
rect 1326 556 1360 590
rect 1484 556 1518 590
rect 1642 556 1676 590
rect 1800 556 1834 590
rect 1958 556 1992 590
rect 2116 556 2150 590
rect 2274 556 2308 590
rect 2432 556 2466 590
rect 2590 556 2624 590
rect 2748 556 2782 590
rect 2906 556 2940 590
rect 3064 556 3098 590
rect -3098 246 -3064 280
rect -2940 246 -2906 280
rect -2782 246 -2748 280
rect -2624 246 -2590 280
rect -2466 246 -2432 280
rect -2308 246 -2274 280
rect -2150 246 -2116 280
rect -1992 246 -1958 280
rect -1834 246 -1800 280
rect -1676 246 -1642 280
rect -1518 246 -1484 280
rect -1360 246 -1326 280
rect -1202 246 -1168 280
rect -1044 246 -1010 280
rect -886 246 -852 280
rect -728 246 -694 280
rect -570 246 -536 280
rect -412 246 -378 280
rect -254 246 -220 280
rect -96 246 -62 280
rect 62 246 96 280
rect 220 246 254 280
rect 378 246 412 280
rect 536 246 570 280
rect 694 246 728 280
rect 852 246 886 280
rect 1010 246 1044 280
rect 1168 246 1202 280
rect 1326 246 1360 280
rect 1484 246 1518 280
rect 1642 246 1676 280
rect 1800 246 1834 280
rect 1958 246 1992 280
rect 2116 246 2150 280
rect 2274 246 2308 280
rect 2432 246 2466 280
rect 2590 246 2624 280
rect 2748 246 2782 280
rect 2906 246 2940 280
rect 3064 246 3098 280
rect -3098 138 -3064 172
rect -2940 138 -2906 172
rect -2782 138 -2748 172
rect -2624 138 -2590 172
rect -2466 138 -2432 172
rect -2308 138 -2274 172
rect -2150 138 -2116 172
rect -1992 138 -1958 172
rect -1834 138 -1800 172
rect -1676 138 -1642 172
rect -1518 138 -1484 172
rect -1360 138 -1326 172
rect -1202 138 -1168 172
rect -1044 138 -1010 172
rect -886 138 -852 172
rect -728 138 -694 172
rect -570 138 -536 172
rect -412 138 -378 172
rect -254 138 -220 172
rect -96 138 -62 172
rect 62 138 96 172
rect 220 138 254 172
rect 378 138 412 172
rect 536 138 570 172
rect 694 138 728 172
rect 852 138 886 172
rect 1010 138 1044 172
rect 1168 138 1202 172
rect 1326 138 1360 172
rect 1484 138 1518 172
rect 1642 138 1676 172
rect 1800 138 1834 172
rect 1958 138 1992 172
rect 2116 138 2150 172
rect 2274 138 2308 172
rect 2432 138 2466 172
rect 2590 138 2624 172
rect 2748 138 2782 172
rect 2906 138 2940 172
rect 3064 138 3098 172
rect -3098 -172 -3064 -138
rect -2940 -172 -2906 -138
rect -2782 -172 -2748 -138
rect -2624 -172 -2590 -138
rect -2466 -172 -2432 -138
rect -2308 -172 -2274 -138
rect -2150 -172 -2116 -138
rect -1992 -172 -1958 -138
rect -1834 -172 -1800 -138
rect -1676 -172 -1642 -138
rect -1518 -172 -1484 -138
rect -1360 -172 -1326 -138
rect -1202 -172 -1168 -138
rect -1044 -172 -1010 -138
rect -886 -172 -852 -138
rect -728 -172 -694 -138
rect -570 -172 -536 -138
rect -412 -172 -378 -138
rect -254 -172 -220 -138
rect -96 -172 -62 -138
rect 62 -172 96 -138
rect 220 -172 254 -138
rect 378 -172 412 -138
rect 536 -172 570 -138
rect 694 -172 728 -138
rect 852 -172 886 -138
rect 1010 -172 1044 -138
rect 1168 -172 1202 -138
rect 1326 -172 1360 -138
rect 1484 -172 1518 -138
rect 1642 -172 1676 -138
rect 1800 -172 1834 -138
rect 1958 -172 1992 -138
rect 2116 -172 2150 -138
rect 2274 -172 2308 -138
rect 2432 -172 2466 -138
rect 2590 -172 2624 -138
rect 2748 -172 2782 -138
rect 2906 -172 2940 -138
rect 3064 -172 3098 -138
rect -3098 -280 -3064 -246
rect -2940 -280 -2906 -246
rect -2782 -280 -2748 -246
rect -2624 -280 -2590 -246
rect -2466 -280 -2432 -246
rect -2308 -280 -2274 -246
rect -2150 -280 -2116 -246
rect -1992 -280 -1958 -246
rect -1834 -280 -1800 -246
rect -1676 -280 -1642 -246
rect -1518 -280 -1484 -246
rect -1360 -280 -1326 -246
rect -1202 -280 -1168 -246
rect -1044 -280 -1010 -246
rect -886 -280 -852 -246
rect -728 -280 -694 -246
rect -570 -280 -536 -246
rect -412 -280 -378 -246
rect -254 -280 -220 -246
rect -96 -280 -62 -246
rect 62 -280 96 -246
rect 220 -280 254 -246
rect 378 -280 412 -246
rect 536 -280 570 -246
rect 694 -280 728 -246
rect 852 -280 886 -246
rect 1010 -280 1044 -246
rect 1168 -280 1202 -246
rect 1326 -280 1360 -246
rect 1484 -280 1518 -246
rect 1642 -280 1676 -246
rect 1800 -280 1834 -246
rect 1958 -280 1992 -246
rect 2116 -280 2150 -246
rect 2274 -280 2308 -246
rect 2432 -280 2466 -246
rect 2590 -280 2624 -246
rect 2748 -280 2782 -246
rect 2906 -280 2940 -246
rect 3064 -280 3098 -246
rect -3098 -590 -3064 -556
rect -2940 -590 -2906 -556
rect -2782 -590 -2748 -556
rect -2624 -590 -2590 -556
rect -2466 -590 -2432 -556
rect -2308 -590 -2274 -556
rect -2150 -590 -2116 -556
rect -1992 -590 -1958 -556
rect -1834 -590 -1800 -556
rect -1676 -590 -1642 -556
rect -1518 -590 -1484 -556
rect -1360 -590 -1326 -556
rect -1202 -590 -1168 -556
rect -1044 -590 -1010 -556
rect -886 -590 -852 -556
rect -728 -590 -694 -556
rect -570 -590 -536 -556
rect -412 -590 -378 -556
rect -254 -590 -220 -556
rect -96 -590 -62 -556
rect 62 -590 96 -556
rect 220 -590 254 -556
rect 378 -590 412 -556
rect 536 -590 570 -556
rect 694 -590 728 -556
rect 852 -590 886 -556
rect 1010 -590 1044 -556
rect 1168 -590 1202 -556
rect 1326 -590 1360 -556
rect 1484 -590 1518 -556
rect 1642 -590 1676 -556
rect 1800 -590 1834 -556
rect 1958 -590 1992 -556
rect 2116 -590 2150 -556
rect 2274 -590 2308 -556
rect 2432 -590 2466 -556
rect 2590 -590 2624 -556
rect 2748 -590 2782 -556
rect 2906 -590 2940 -556
rect 3064 -590 3098 -556
<< locali >>
rect -3311 694 -3213 728
rect -3179 694 -3145 728
rect -3111 694 -3077 728
rect -3043 694 -3009 728
rect -2975 694 -2941 728
rect -2907 694 -2873 728
rect -2839 694 -2805 728
rect -2771 694 -2737 728
rect -2703 694 -2669 728
rect -2635 694 -2601 728
rect -2567 694 -2533 728
rect -2499 694 -2465 728
rect -2431 694 -2397 728
rect -2363 694 -2329 728
rect -2295 694 -2261 728
rect -2227 694 -2193 728
rect -2159 694 -2125 728
rect -2091 694 -2057 728
rect -2023 694 -1989 728
rect -1955 694 -1921 728
rect -1887 694 -1853 728
rect -1819 694 -1785 728
rect -1751 694 -1717 728
rect -1683 694 -1649 728
rect -1615 694 -1581 728
rect -1547 694 -1513 728
rect -1479 694 -1445 728
rect -1411 694 -1377 728
rect -1343 694 -1309 728
rect -1275 694 -1241 728
rect -1207 694 -1173 728
rect -1139 694 -1105 728
rect -1071 694 -1037 728
rect -1003 694 -969 728
rect -935 694 -901 728
rect -867 694 -833 728
rect -799 694 -765 728
rect -731 694 -697 728
rect -663 694 -629 728
rect -595 694 -561 728
rect -527 694 -493 728
rect -459 694 -425 728
rect -391 694 -357 728
rect -323 694 -289 728
rect -255 694 -221 728
rect -187 694 -153 728
rect -119 694 -85 728
rect -51 694 -17 728
rect 17 694 51 728
rect 85 694 119 728
rect 153 694 187 728
rect 221 694 255 728
rect 289 694 323 728
rect 357 694 391 728
rect 425 694 459 728
rect 493 694 527 728
rect 561 694 595 728
rect 629 694 663 728
rect 697 694 731 728
rect 765 694 799 728
rect 833 694 867 728
rect 901 694 935 728
rect 969 694 1003 728
rect 1037 694 1071 728
rect 1105 694 1139 728
rect 1173 694 1207 728
rect 1241 694 1275 728
rect 1309 694 1343 728
rect 1377 694 1411 728
rect 1445 694 1479 728
rect 1513 694 1547 728
rect 1581 694 1615 728
rect 1649 694 1683 728
rect 1717 694 1751 728
rect 1785 694 1819 728
rect 1853 694 1887 728
rect 1921 694 1955 728
rect 1989 694 2023 728
rect 2057 694 2091 728
rect 2125 694 2159 728
rect 2193 694 2227 728
rect 2261 694 2295 728
rect 2329 694 2363 728
rect 2397 694 2431 728
rect 2465 694 2499 728
rect 2533 694 2567 728
rect 2601 694 2635 728
rect 2669 694 2703 728
rect 2737 694 2771 728
rect 2805 694 2839 728
rect 2873 694 2907 728
rect 2941 694 2975 728
rect 3009 694 3043 728
rect 3077 694 3111 728
rect 3145 694 3179 728
rect 3213 694 3311 728
rect -3311 629 -3277 694
rect -3311 561 -3277 595
rect 3277 629 3311 694
rect -3131 556 -3098 590
rect -3064 556 -3031 590
rect -2973 556 -2940 590
rect -2906 556 -2873 590
rect -2815 556 -2782 590
rect -2748 556 -2715 590
rect -2657 556 -2624 590
rect -2590 556 -2557 590
rect -2499 556 -2466 590
rect -2432 556 -2399 590
rect -2341 556 -2308 590
rect -2274 556 -2241 590
rect -2183 556 -2150 590
rect -2116 556 -2083 590
rect -2025 556 -1992 590
rect -1958 556 -1925 590
rect -1867 556 -1834 590
rect -1800 556 -1767 590
rect -1709 556 -1676 590
rect -1642 556 -1609 590
rect -1551 556 -1518 590
rect -1484 556 -1451 590
rect -1393 556 -1360 590
rect -1326 556 -1293 590
rect -1235 556 -1202 590
rect -1168 556 -1135 590
rect -1077 556 -1044 590
rect -1010 556 -977 590
rect -919 556 -886 590
rect -852 556 -819 590
rect -761 556 -728 590
rect -694 556 -661 590
rect -603 556 -570 590
rect -536 556 -503 590
rect -445 556 -412 590
rect -378 556 -345 590
rect -287 556 -254 590
rect -220 556 -187 590
rect -129 556 -96 590
rect -62 556 -29 590
rect 29 556 62 590
rect 96 556 129 590
rect 187 556 220 590
rect 254 556 287 590
rect 345 556 378 590
rect 412 556 445 590
rect 503 556 536 590
rect 570 556 603 590
rect 661 556 694 590
rect 728 556 761 590
rect 819 556 852 590
rect 886 556 919 590
rect 977 556 1010 590
rect 1044 556 1077 590
rect 1135 556 1168 590
rect 1202 556 1235 590
rect 1293 556 1326 590
rect 1360 556 1393 590
rect 1451 556 1484 590
rect 1518 556 1551 590
rect 1609 556 1642 590
rect 1676 556 1709 590
rect 1767 556 1800 590
rect 1834 556 1867 590
rect 1925 556 1958 590
rect 1992 556 2025 590
rect 2083 556 2116 590
rect 2150 556 2183 590
rect 2241 556 2274 590
rect 2308 556 2341 590
rect 2399 556 2432 590
rect 2466 556 2499 590
rect 2557 556 2590 590
rect 2624 556 2657 590
rect 2715 556 2748 590
rect 2782 556 2815 590
rect 2873 556 2906 590
rect 2940 556 2973 590
rect 3031 556 3064 590
rect 3098 556 3131 590
rect 3277 561 3311 595
rect -3311 493 -3277 527
rect -3311 425 -3277 459
rect -3311 357 -3277 391
rect -3311 289 -3277 323
rect -3177 503 -3143 522
rect -3177 435 -3143 437
rect -3177 399 -3143 401
rect -3177 314 -3143 333
rect -3019 503 -2985 522
rect -3019 435 -2985 437
rect -3019 399 -2985 401
rect -3019 314 -2985 333
rect -2861 503 -2827 522
rect -2861 435 -2827 437
rect -2861 399 -2827 401
rect -2861 314 -2827 333
rect -2703 503 -2669 522
rect -2703 435 -2669 437
rect -2703 399 -2669 401
rect -2703 314 -2669 333
rect -2545 503 -2511 522
rect -2545 435 -2511 437
rect -2545 399 -2511 401
rect -2545 314 -2511 333
rect -2387 503 -2353 522
rect -2387 435 -2353 437
rect -2387 399 -2353 401
rect -2387 314 -2353 333
rect -2229 503 -2195 522
rect -2229 435 -2195 437
rect -2229 399 -2195 401
rect -2229 314 -2195 333
rect -2071 503 -2037 522
rect -2071 435 -2037 437
rect -2071 399 -2037 401
rect -2071 314 -2037 333
rect -1913 503 -1879 522
rect -1913 435 -1879 437
rect -1913 399 -1879 401
rect -1913 314 -1879 333
rect -1755 503 -1721 522
rect -1755 435 -1721 437
rect -1755 399 -1721 401
rect -1755 314 -1721 333
rect -1597 503 -1563 522
rect -1597 435 -1563 437
rect -1597 399 -1563 401
rect -1597 314 -1563 333
rect -1439 503 -1405 522
rect -1439 435 -1405 437
rect -1439 399 -1405 401
rect -1439 314 -1405 333
rect -1281 503 -1247 522
rect -1281 435 -1247 437
rect -1281 399 -1247 401
rect -1281 314 -1247 333
rect -1123 503 -1089 522
rect -1123 435 -1089 437
rect -1123 399 -1089 401
rect -1123 314 -1089 333
rect -965 503 -931 522
rect -965 435 -931 437
rect -965 399 -931 401
rect -965 314 -931 333
rect -807 503 -773 522
rect -807 435 -773 437
rect -807 399 -773 401
rect -807 314 -773 333
rect -649 503 -615 522
rect -649 435 -615 437
rect -649 399 -615 401
rect -649 314 -615 333
rect -491 503 -457 522
rect -491 435 -457 437
rect -491 399 -457 401
rect -491 314 -457 333
rect -333 503 -299 522
rect -333 435 -299 437
rect -333 399 -299 401
rect -333 314 -299 333
rect -175 503 -141 522
rect -175 435 -141 437
rect -175 399 -141 401
rect -175 314 -141 333
rect -17 503 17 522
rect -17 435 17 437
rect -17 399 17 401
rect -17 314 17 333
rect 141 503 175 522
rect 141 435 175 437
rect 141 399 175 401
rect 141 314 175 333
rect 299 503 333 522
rect 299 435 333 437
rect 299 399 333 401
rect 299 314 333 333
rect 457 503 491 522
rect 457 435 491 437
rect 457 399 491 401
rect 457 314 491 333
rect 615 503 649 522
rect 615 435 649 437
rect 615 399 649 401
rect 615 314 649 333
rect 773 503 807 522
rect 773 435 807 437
rect 773 399 807 401
rect 773 314 807 333
rect 931 503 965 522
rect 931 435 965 437
rect 931 399 965 401
rect 931 314 965 333
rect 1089 503 1123 522
rect 1089 435 1123 437
rect 1089 399 1123 401
rect 1089 314 1123 333
rect 1247 503 1281 522
rect 1247 435 1281 437
rect 1247 399 1281 401
rect 1247 314 1281 333
rect 1405 503 1439 522
rect 1405 435 1439 437
rect 1405 399 1439 401
rect 1405 314 1439 333
rect 1563 503 1597 522
rect 1563 435 1597 437
rect 1563 399 1597 401
rect 1563 314 1597 333
rect 1721 503 1755 522
rect 1721 435 1755 437
rect 1721 399 1755 401
rect 1721 314 1755 333
rect 1879 503 1913 522
rect 1879 435 1913 437
rect 1879 399 1913 401
rect 1879 314 1913 333
rect 2037 503 2071 522
rect 2037 435 2071 437
rect 2037 399 2071 401
rect 2037 314 2071 333
rect 2195 503 2229 522
rect 2195 435 2229 437
rect 2195 399 2229 401
rect 2195 314 2229 333
rect 2353 503 2387 522
rect 2353 435 2387 437
rect 2353 399 2387 401
rect 2353 314 2387 333
rect 2511 503 2545 522
rect 2511 435 2545 437
rect 2511 399 2545 401
rect 2511 314 2545 333
rect 2669 503 2703 522
rect 2669 435 2703 437
rect 2669 399 2703 401
rect 2669 314 2703 333
rect 2827 503 2861 522
rect 2827 435 2861 437
rect 2827 399 2861 401
rect 2827 314 2861 333
rect 2985 503 3019 522
rect 2985 435 3019 437
rect 2985 399 3019 401
rect 2985 314 3019 333
rect 3143 503 3177 522
rect 3143 435 3177 437
rect 3143 399 3177 401
rect 3143 314 3177 333
rect 3277 493 3311 527
rect 3277 425 3311 459
rect 3277 357 3311 391
rect 3277 289 3311 323
rect -3311 221 -3277 255
rect -3131 246 -3098 280
rect -3064 246 -3031 280
rect -2973 246 -2940 280
rect -2906 246 -2873 280
rect -2815 246 -2782 280
rect -2748 246 -2715 280
rect -2657 246 -2624 280
rect -2590 246 -2557 280
rect -2499 246 -2466 280
rect -2432 246 -2399 280
rect -2341 246 -2308 280
rect -2274 246 -2241 280
rect -2183 246 -2150 280
rect -2116 246 -2083 280
rect -2025 246 -1992 280
rect -1958 246 -1925 280
rect -1867 246 -1834 280
rect -1800 246 -1767 280
rect -1709 246 -1676 280
rect -1642 246 -1609 280
rect -1551 246 -1518 280
rect -1484 246 -1451 280
rect -1393 246 -1360 280
rect -1326 246 -1293 280
rect -1235 246 -1202 280
rect -1168 246 -1135 280
rect -1077 246 -1044 280
rect -1010 246 -977 280
rect -919 246 -886 280
rect -852 246 -819 280
rect -761 246 -728 280
rect -694 246 -661 280
rect -603 246 -570 280
rect -536 246 -503 280
rect -445 246 -412 280
rect -378 246 -345 280
rect -287 246 -254 280
rect -220 246 -187 280
rect -129 246 -96 280
rect -62 246 -29 280
rect 29 246 62 280
rect 96 246 129 280
rect 187 246 220 280
rect 254 246 287 280
rect 345 246 378 280
rect 412 246 445 280
rect 503 246 536 280
rect 570 246 603 280
rect 661 246 694 280
rect 728 246 761 280
rect 819 246 852 280
rect 886 246 919 280
rect 977 246 1010 280
rect 1044 246 1077 280
rect 1135 246 1168 280
rect 1202 246 1235 280
rect 1293 246 1326 280
rect 1360 246 1393 280
rect 1451 246 1484 280
rect 1518 246 1551 280
rect 1609 246 1642 280
rect 1676 246 1709 280
rect 1767 246 1800 280
rect 1834 246 1867 280
rect 1925 246 1958 280
rect 1992 246 2025 280
rect 2083 246 2116 280
rect 2150 246 2183 280
rect 2241 246 2274 280
rect 2308 246 2341 280
rect 2399 246 2432 280
rect 2466 246 2499 280
rect 2557 246 2590 280
rect 2624 246 2657 280
rect 2715 246 2748 280
rect 2782 246 2815 280
rect 2873 246 2906 280
rect 2940 246 2973 280
rect 3031 246 3064 280
rect 3098 246 3131 280
rect -3311 153 -3277 187
rect 3277 221 3311 255
rect -3131 138 -3098 172
rect -3064 138 -3031 172
rect -2973 138 -2940 172
rect -2906 138 -2873 172
rect -2815 138 -2782 172
rect -2748 138 -2715 172
rect -2657 138 -2624 172
rect -2590 138 -2557 172
rect -2499 138 -2466 172
rect -2432 138 -2399 172
rect -2341 138 -2308 172
rect -2274 138 -2241 172
rect -2183 138 -2150 172
rect -2116 138 -2083 172
rect -2025 138 -1992 172
rect -1958 138 -1925 172
rect -1867 138 -1834 172
rect -1800 138 -1767 172
rect -1709 138 -1676 172
rect -1642 138 -1609 172
rect -1551 138 -1518 172
rect -1484 138 -1451 172
rect -1393 138 -1360 172
rect -1326 138 -1293 172
rect -1235 138 -1202 172
rect -1168 138 -1135 172
rect -1077 138 -1044 172
rect -1010 138 -977 172
rect -919 138 -886 172
rect -852 138 -819 172
rect -761 138 -728 172
rect -694 138 -661 172
rect -603 138 -570 172
rect -536 138 -503 172
rect -445 138 -412 172
rect -378 138 -345 172
rect -287 138 -254 172
rect -220 138 -187 172
rect -129 138 -96 172
rect -62 138 -29 172
rect 29 138 62 172
rect 96 138 129 172
rect 187 138 220 172
rect 254 138 287 172
rect 345 138 378 172
rect 412 138 445 172
rect 503 138 536 172
rect 570 138 603 172
rect 661 138 694 172
rect 728 138 761 172
rect 819 138 852 172
rect 886 138 919 172
rect 977 138 1010 172
rect 1044 138 1077 172
rect 1135 138 1168 172
rect 1202 138 1235 172
rect 1293 138 1326 172
rect 1360 138 1393 172
rect 1451 138 1484 172
rect 1518 138 1551 172
rect 1609 138 1642 172
rect 1676 138 1709 172
rect 1767 138 1800 172
rect 1834 138 1867 172
rect 1925 138 1958 172
rect 1992 138 2025 172
rect 2083 138 2116 172
rect 2150 138 2183 172
rect 2241 138 2274 172
rect 2308 138 2341 172
rect 2399 138 2432 172
rect 2466 138 2499 172
rect 2557 138 2590 172
rect 2624 138 2657 172
rect 2715 138 2748 172
rect 2782 138 2815 172
rect 2873 138 2906 172
rect 2940 138 2973 172
rect 3031 138 3064 172
rect 3098 138 3131 172
rect 3277 153 3311 187
rect -3311 85 -3277 119
rect -3311 17 -3277 51
rect -3311 -51 -3277 -17
rect -3311 -119 -3277 -85
rect -3177 85 -3143 104
rect -3177 17 -3143 19
rect -3177 -19 -3143 -17
rect -3177 -104 -3143 -85
rect -3019 85 -2985 104
rect -3019 17 -2985 19
rect -3019 -19 -2985 -17
rect -3019 -104 -2985 -85
rect -2861 85 -2827 104
rect -2861 17 -2827 19
rect -2861 -19 -2827 -17
rect -2861 -104 -2827 -85
rect -2703 85 -2669 104
rect -2703 17 -2669 19
rect -2703 -19 -2669 -17
rect -2703 -104 -2669 -85
rect -2545 85 -2511 104
rect -2545 17 -2511 19
rect -2545 -19 -2511 -17
rect -2545 -104 -2511 -85
rect -2387 85 -2353 104
rect -2387 17 -2353 19
rect -2387 -19 -2353 -17
rect -2387 -104 -2353 -85
rect -2229 85 -2195 104
rect -2229 17 -2195 19
rect -2229 -19 -2195 -17
rect -2229 -104 -2195 -85
rect -2071 85 -2037 104
rect -2071 17 -2037 19
rect -2071 -19 -2037 -17
rect -2071 -104 -2037 -85
rect -1913 85 -1879 104
rect -1913 17 -1879 19
rect -1913 -19 -1879 -17
rect -1913 -104 -1879 -85
rect -1755 85 -1721 104
rect -1755 17 -1721 19
rect -1755 -19 -1721 -17
rect -1755 -104 -1721 -85
rect -1597 85 -1563 104
rect -1597 17 -1563 19
rect -1597 -19 -1563 -17
rect -1597 -104 -1563 -85
rect -1439 85 -1405 104
rect -1439 17 -1405 19
rect -1439 -19 -1405 -17
rect -1439 -104 -1405 -85
rect -1281 85 -1247 104
rect -1281 17 -1247 19
rect -1281 -19 -1247 -17
rect -1281 -104 -1247 -85
rect -1123 85 -1089 104
rect -1123 17 -1089 19
rect -1123 -19 -1089 -17
rect -1123 -104 -1089 -85
rect -965 85 -931 104
rect -965 17 -931 19
rect -965 -19 -931 -17
rect -965 -104 -931 -85
rect -807 85 -773 104
rect -807 17 -773 19
rect -807 -19 -773 -17
rect -807 -104 -773 -85
rect -649 85 -615 104
rect -649 17 -615 19
rect -649 -19 -615 -17
rect -649 -104 -615 -85
rect -491 85 -457 104
rect -491 17 -457 19
rect -491 -19 -457 -17
rect -491 -104 -457 -85
rect -333 85 -299 104
rect -333 17 -299 19
rect -333 -19 -299 -17
rect -333 -104 -299 -85
rect -175 85 -141 104
rect -175 17 -141 19
rect -175 -19 -141 -17
rect -175 -104 -141 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 141 85 175 104
rect 141 17 175 19
rect 141 -19 175 -17
rect 141 -104 175 -85
rect 299 85 333 104
rect 299 17 333 19
rect 299 -19 333 -17
rect 299 -104 333 -85
rect 457 85 491 104
rect 457 17 491 19
rect 457 -19 491 -17
rect 457 -104 491 -85
rect 615 85 649 104
rect 615 17 649 19
rect 615 -19 649 -17
rect 615 -104 649 -85
rect 773 85 807 104
rect 773 17 807 19
rect 773 -19 807 -17
rect 773 -104 807 -85
rect 931 85 965 104
rect 931 17 965 19
rect 931 -19 965 -17
rect 931 -104 965 -85
rect 1089 85 1123 104
rect 1089 17 1123 19
rect 1089 -19 1123 -17
rect 1089 -104 1123 -85
rect 1247 85 1281 104
rect 1247 17 1281 19
rect 1247 -19 1281 -17
rect 1247 -104 1281 -85
rect 1405 85 1439 104
rect 1405 17 1439 19
rect 1405 -19 1439 -17
rect 1405 -104 1439 -85
rect 1563 85 1597 104
rect 1563 17 1597 19
rect 1563 -19 1597 -17
rect 1563 -104 1597 -85
rect 1721 85 1755 104
rect 1721 17 1755 19
rect 1721 -19 1755 -17
rect 1721 -104 1755 -85
rect 1879 85 1913 104
rect 1879 17 1913 19
rect 1879 -19 1913 -17
rect 1879 -104 1913 -85
rect 2037 85 2071 104
rect 2037 17 2071 19
rect 2037 -19 2071 -17
rect 2037 -104 2071 -85
rect 2195 85 2229 104
rect 2195 17 2229 19
rect 2195 -19 2229 -17
rect 2195 -104 2229 -85
rect 2353 85 2387 104
rect 2353 17 2387 19
rect 2353 -19 2387 -17
rect 2353 -104 2387 -85
rect 2511 85 2545 104
rect 2511 17 2545 19
rect 2511 -19 2545 -17
rect 2511 -104 2545 -85
rect 2669 85 2703 104
rect 2669 17 2703 19
rect 2669 -19 2703 -17
rect 2669 -104 2703 -85
rect 2827 85 2861 104
rect 2827 17 2861 19
rect 2827 -19 2861 -17
rect 2827 -104 2861 -85
rect 2985 85 3019 104
rect 2985 17 3019 19
rect 2985 -19 3019 -17
rect 2985 -104 3019 -85
rect 3143 85 3177 104
rect 3143 17 3177 19
rect 3143 -19 3177 -17
rect 3143 -104 3177 -85
rect 3277 85 3311 119
rect 3277 17 3311 51
rect 3277 -51 3311 -17
rect 3277 -119 3311 -85
rect -3311 -187 -3277 -153
rect -3131 -172 -3098 -138
rect -3064 -172 -3031 -138
rect -2973 -172 -2940 -138
rect -2906 -172 -2873 -138
rect -2815 -172 -2782 -138
rect -2748 -172 -2715 -138
rect -2657 -172 -2624 -138
rect -2590 -172 -2557 -138
rect -2499 -172 -2466 -138
rect -2432 -172 -2399 -138
rect -2341 -172 -2308 -138
rect -2274 -172 -2241 -138
rect -2183 -172 -2150 -138
rect -2116 -172 -2083 -138
rect -2025 -172 -1992 -138
rect -1958 -172 -1925 -138
rect -1867 -172 -1834 -138
rect -1800 -172 -1767 -138
rect -1709 -172 -1676 -138
rect -1642 -172 -1609 -138
rect -1551 -172 -1518 -138
rect -1484 -172 -1451 -138
rect -1393 -172 -1360 -138
rect -1326 -172 -1293 -138
rect -1235 -172 -1202 -138
rect -1168 -172 -1135 -138
rect -1077 -172 -1044 -138
rect -1010 -172 -977 -138
rect -919 -172 -886 -138
rect -852 -172 -819 -138
rect -761 -172 -728 -138
rect -694 -172 -661 -138
rect -603 -172 -570 -138
rect -536 -172 -503 -138
rect -445 -172 -412 -138
rect -378 -172 -345 -138
rect -287 -172 -254 -138
rect -220 -172 -187 -138
rect -129 -172 -96 -138
rect -62 -172 -29 -138
rect 29 -172 62 -138
rect 96 -172 129 -138
rect 187 -172 220 -138
rect 254 -172 287 -138
rect 345 -172 378 -138
rect 412 -172 445 -138
rect 503 -172 536 -138
rect 570 -172 603 -138
rect 661 -172 694 -138
rect 728 -172 761 -138
rect 819 -172 852 -138
rect 886 -172 919 -138
rect 977 -172 1010 -138
rect 1044 -172 1077 -138
rect 1135 -172 1168 -138
rect 1202 -172 1235 -138
rect 1293 -172 1326 -138
rect 1360 -172 1393 -138
rect 1451 -172 1484 -138
rect 1518 -172 1551 -138
rect 1609 -172 1642 -138
rect 1676 -172 1709 -138
rect 1767 -172 1800 -138
rect 1834 -172 1867 -138
rect 1925 -172 1958 -138
rect 1992 -172 2025 -138
rect 2083 -172 2116 -138
rect 2150 -172 2183 -138
rect 2241 -172 2274 -138
rect 2308 -172 2341 -138
rect 2399 -172 2432 -138
rect 2466 -172 2499 -138
rect 2557 -172 2590 -138
rect 2624 -172 2657 -138
rect 2715 -172 2748 -138
rect 2782 -172 2815 -138
rect 2873 -172 2906 -138
rect 2940 -172 2973 -138
rect 3031 -172 3064 -138
rect 3098 -172 3131 -138
rect -3311 -255 -3277 -221
rect 3277 -187 3311 -153
rect -3131 -280 -3098 -246
rect -3064 -280 -3031 -246
rect -2973 -280 -2940 -246
rect -2906 -280 -2873 -246
rect -2815 -280 -2782 -246
rect -2748 -280 -2715 -246
rect -2657 -280 -2624 -246
rect -2590 -280 -2557 -246
rect -2499 -280 -2466 -246
rect -2432 -280 -2399 -246
rect -2341 -280 -2308 -246
rect -2274 -280 -2241 -246
rect -2183 -280 -2150 -246
rect -2116 -280 -2083 -246
rect -2025 -280 -1992 -246
rect -1958 -280 -1925 -246
rect -1867 -280 -1834 -246
rect -1800 -280 -1767 -246
rect -1709 -280 -1676 -246
rect -1642 -280 -1609 -246
rect -1551 -280 -1518 -246
rect -1484 -280 -1451 -246
rect -1393 -280 -1360 -246
rect -1326 -280 -1293 -246
rect -1235 -280 -1202 -246
rect -1168 -280 -1135 -246
rect -1077 -280 -1044 -246
rect -1010 -280 -977 -246
rect -919 -280 -886 -246
rect -852 -280 -819 -246
rect -761 -280 -728 -246
rect -694 -280 -661 -246
rect -603 -280 -570 -246
rect -536 -280 -503 -246
rect -445 -280 -412 -246
rect -378 -280 -345 -246
rect -287 -280 -254 -246
rect -220 -280 -187 -246
rect -129 -280 -96 -246
rect -62 -280 -29 -246
rect 29 -280 62 -246
rect 96 -280 129 -246
rect 187 -280 220 -246
rect 254 -280 287 -246
rect 345 -280 378 -246
rect 412 -280 445 -246
rect 503 -280 536 -246
rect 570 -280 603 -246
rect 661 -280 694 -246
rect 728 -280 761 -246
rect 819 -280 852 -246
rect 886 -280 919 -246
rect 977 -280 1010 -246
rect 1044 -280 1077 -246
rect 1135 -280 1168 -246
rect 1202 -280 1235 -246
rect 1293 -280 1326 -246
rect 1360 -280 1393 -246
rect 1451 -280 1484 -246
rect 1518 -280 1551 -246
rect 1609 -280 1642 -246
rect 1676 -280 1709 -246
rect 1767 -280 1800 -246
rect 1834 -280 1867 -246
rect 1925 -280 1958 -246
rect 1992 -280 2025 -246
rect 2083 -280 2116 -246
rect 2150 -280 2183 -246
rect 2241 -280 2274 -246
rect 2308 -280 2341 -246
rect 2399 -280 2432 -246
rect 2466 -280 2499 -246
rect 2557 -280 2590 -246
rect 2624 -280 2657 -246
rect 2715 -280 2748 -246
rect 2782 -280 2815 -246
rect 2873 -280 2906 -246
rect 2940 -280 2973 -246
rect 3031 -280 3064 -246
rect 3098 -280 3131 -246
rect 3277 -255 3311 -221
rect -3311 -323 -3277 -289
rect -3311 -391 -3277 -357
rect -3311 -459 -3277 -425
rect -3311 -527 -3277 -493
rect -3177 -333 -3143 -314
rect -3177 -401 -3143 -399
rect -3177 -437 -3143 -435
rect -3177 -522 -3143 -503
rect -3019 -333 -2985 -314
rect -3019 -401 -2985 -399
rect -3019 -437 -2985 -435
rect -3019 -522 -2985 -503
rect -2861 -333 -2827 -314
rect -2861 -401 -2827 -399
rect -2861 -437 -2827 -435
rect -2861 -522 -2827 -503
rect -2703 -333 -2669 -314
rect -2703 -401 -2669 -399
rect -2703 -437 -2669 -435
rect -2703 -522 -2669 -503
rect -2545 -333 -2511 -314
rect -2545 -401 -2511 -399
rect -2545 -437 -2511 -435
rect -2545 -522 -2511 -503
rect -2387 -333 -2353 -314
rect -2387 -401 -2353 -399
rect -2387 -437 -2353 -435
rect -2387 -522 -2353 -503
rect -2229 -333 -2195 -314
rect -2229 -401 -2195 -399
rect -2229 -437 -2195 -435
rect -2229 -522 -2195 -503
rect -2071 -333 -2037 -314
rect -2071 -401 -2037 -399
rect -2071 -437 -2037 -435
rect -2071 -522 -2037 -503
rect -1913 -333 -1879 -314
rect -1913 -401 -1879 -399
rect -1913 -437 -1879 -435
rect -1913 -522 -1879 -503
rect -1755 -333 -1721 -314
rect -1755 -401 -1721 -399
rect -1755 -437 -1721 -435
rect -1755 -522 -1721 -503
rect -1597 -333 -1563 -314
rect -1597 -401 -1563 -399
rect -1597 -437 -1563 -435
rect -1597 -522 -1563 -503
rect -1439 -333 -1405 -314
rect -1439 -401 -1405 -399
rect -1439 -437 -1405 -435
rect -1439 -522 -1405 -503
rect -1281 -333 -1247 -314
rect -1281 -401 -1247 -399
rect -1281 -437 -1247 -435
rect -1281 -522 -1247 -503
rect -1123 -333 -1089 -314
rect -1123 -401 -1089 -399
rect -1123 -437 -1089 -435
rect -1123 -522 -1089 -503
rect -965 -333 -931 -314
rect -965 -401 -931 -399
rect -965 -437 -931 -435
rect -965 -522 -931 -503
rect -807 -333 -773 -314
rect -807 -401 -773 -399
rect -807 -437 -773 -435
rect -807 -522 -773 -503
rect -649 -333 -615 -314
rect -649 -401 -615 -399
rect -649 -437 -615 -435
rect -649 -522 -615 -503
rect -491 -333 -457 -314
rect -491 -401 -457 -399
rect -491 -437 -457 -435
rect -491 -522 -457 -503
rect -333 -333 -299 -314
rect -333 -401 -299 -399
rect -333 -437 -299 -435
rect -333 -522 -299 -503
rect -175 -333 -141 -314
rect -175 -401 -141 -399
rect -175 -437 -141 -435
rect -175 -522 -141 -503
rect -17 -333 17 -314
rect -17 -401 17 -399
rect -17 -437 17 -435
rect -17 -522 17 -503
rect 141 -333 175 -314
rect 141 -401 175 -399
rect 141 -437 175 -435
rect 141 -522 175 -503
rect 299 -333 333 -314
rect 299 -401 333 -399
rect 299 -437 333 -435
rect 299 -522 333 -503
rect 457 -333 491 -314
rect 457 -401 491 -399
rect 457 -437 491 -435
rect 457 -522 491 -503
rect 615 -333 649 -314
rect 615 -401 649 -399
rect 615 -437 649 -435
rect 615 -522 649 -503
rect 773 -333 807 -314
rect 773 -401 807 -399
rect 773 -437 807 -435
rect 773 -522 807 -503
rect 931 -333 965 -314
rect 931 -401 965 -399
rect 931 -437 965 -435
rect 931 -522 965 -503
rect 1089 -333 1123 -314
rect 1089 -401 1123 -399
rect 1089 -437 1123 -435
rect 1089 -522 1123 -503
rect 1247 -333 1281 -314
rect 1247 -401 1281 -399
rect 1247 -437 1281 -435
rect 1247 -522 1281 -503
rect 1405 -333 1439 -314
rect 1405 -401 1439 -399
rect 1405 -437 1439 -435
rect 1405 -522 1439 -503
rect 1563 -333 1597 -314
rect 1563 -401 1597 -399
rect 1563 -437 1597 -435
rect 1563 -522 1597 -503
rect 1721 -333 1755 -314
rect 1721 -401 1755 -399
rect 1721 -437 1755 -435
rect 1721 -522 1755 -503
rect 1879 -333 1913 -314
rect 1879 -401 1913 -399
rect 1879 -437 1913 -435
rect 1879 -522 1913 -503
rect 2037 -333 2071 -314
rect 2037 -401 2071 -399
rect 2037 -437 2071 -435
rect 2037 -522 2071 -503
rect 2195 -333 2229 -314
rect 2195 -401 2229 -399
rect 2195 -437 2229 -435
rect 2195 -522 2229 -503
rect 2353 -333 2387 -314
rect 2353 -401 2387 -399
rect 2353 -437 2387 -435
rect 2353 -522 2387 -503
rect 2511 -333 2545 -314
rect 2511 -401 2545 -399
rect 2511 -437 2545 -435
rect 2511 -522 2545 -503
rect 2669 -333 2703 -314
rect 2669 -401 2703 -399
rect 2669 -437 2703 -435
rect 2669 -522 2703 -503
rect 2827 -333 2861 -314
rect 2827 -401 2861 -399
rect 2827 -437 2861 -435
rect 2827 -522 2861 -503
rect 2985 -333 3019 -314
rect 2985 -401 3019 -399
rect 2985 -437 3019 -435
rect 2985 -522 3019 -503
rect 3143 -333 3177 -314
rect 3143 -401 3177 -399
rect 3143 -437 3177 -435
rect 3143 -522 3177 -503
rect 3277 -323 3311 -289
rect 3277 -391 3311 -357
rect 3277 -459 3311 -425
rect 3277 -527 3311 -493
rect -3311 -595 -3277 -561
rect -3131 -590 -3098 -556
rect -3064 -590 -3031 -556
rect -2973 -590 -2940 -556
rect -2906 -590 -2873 -556
rect -2815 -590 -2782 -556
rect -2748 -590 -2715 -556
rect -2657 -590 -2624 -556
rect -2590 -590 -2557 -556
rect -2499 -590 -2466 -556
rect -2432 -590 -2399 -556
rect -2341 -590 -2308 -556
rect -2274 -590 -2241 -556
rect -2183 -590 -2150 -556
rect -2116 -590 -2083 -556
rect -2025 -590 -1992 -556
rect -1958 -590 -1925 -556
rect -1867 -590 -1834 -556
rect -1800 -590 -1767 -556
rect -1709 -590 -1676 -556
rect -1642 -590 -1609 -556
rect -1551 -590 -1518 -556
rect -1484 -590 -1451 -556
rect -1393 -590 -1360 -556
rect -1326 -590 -1293 -556
rect -1235 -590 -1202 -556
rect -1168 -590 -1135 -556
rect -1077 -590 -1044 -556
rect -1010 -590 -977 -556
rect -919 -590 -886 -556
rect -852 -590 -819 -556
rect -761 -590 -728 -556
rect -694 -590 -661 -556
rect -603 -590 -570 -556
rect -536 -590 -503 -556
rect -445 -590 -412 -556
rect -378 -590 -345 -556
rect -287 -590 -254 -556
rect -220 -590 -187 -556
rect -129 -590 -96 -556
rect -62 -590 -29 -556
rect 29 -590 62 -556
rect 96 -590 129 -556
rect 187 -590 220 -556
rect 254 -590 287 -556
rect 345 -590 378 -556
rect 412 -590 445 -556
rect 503 -590 536 -556
rect 570 -590 603 -556
rect 661 -590 694 -556
rect 728 -590 761 -556
rect 819 -590 852 -556
rect 886 -590 919 -556
rect 977 -590 1010 -556
rect 1044 -590 1077 -556
rect 1135 -590 1168 -556
rect 1202 -590 1235 -556
rect 1293 -590 1326 -556
rect 1360 -590 1393 -556
rect 1451 -590 1484 -556
rect 1518 -590 1551 -556
rect 1609 -590 1642 -556
rect 1676 -590 1709 -556
rect 1767 -590 1800 -556
rect 1834 -590 1867 -556
rect 1925 -590 1958 -556
rect 1992 -590 2025 -556
rect 2083 -590 2116 -556
rect 2150 -590 2183 -556
rect 2241 -590 2274 -556
rect 2308 -590 2341 -556
rect 2399 -590 2432 -556
rect 2466 -590 2499 -556
rect 2557 -590 2590 -556
rect 2624 -590 2657 -556
rect 2715 -590 2748 -556
rect 2782 -590 2815 -556
rect 2873 -590 2906 -556
rect 2940 -590 2973 -556
rect 3031 -590 3064 -556
rect 3098 -590 3131 -556
rect -3311 -694 -3277 -629
rect 3277 -595 3311 -561
rect 3277 -694 3311 -629
rect -3311 -728 -3213 -694
rect -3179 -728 -3145 -694
rect -3111 -728 -3077 -694
rect -3043 -728 -3009 -694
rect -2975 -728 -2941 -694
rect -2907 -728 -2873 -694
rect -2839 -728 -2805 -694
rect -2771 -728 -2737 -694
rect -2703 -728 -2669 -694
rect -2635 -728 -2601 -694
rect -2567 -728 -2533 -694
rect -2499 -728 -2465 -694
rect -2431 -728 -2397 -694
rect -2363 -728 -2329 -694
rect -2295 -728 -2261 -694
rect -2227 -728 -2193 -694
rect -2159 -728 -2125 -694
rect -2091 -728 -2057 -694
rect -2023 -728 -1989 -694
rect -1955 -728 -1921 -694
rect -1887 -728 -1853 -694
rect -1819 -728 -1785 -694
rect -1751 -728 -1717 -694
rect -1683 -728 -1649 -694
rect -1615 -728 -1581 -694
rect -1547 -728 -1513 -694
rect -1479 -728 -1445 -694
rect -1411 -728 -1377 -694
rect -1343 -728 -1309 -694
rect -1275 -728 -1241 -694
rect -1207 -728 -1173 -694
rect -1139 -728 -1105 -694
rect -1071 -728 -1037 -694
rect -1003 -728 -969 -694
rect -935 -728 -901 -694
rect -867 -728 -833 -694
rect -799 -728 -765 -694
rect -731 -728 -697 -694
rect -663 -728 -629 -694
rect -595 -728 -561 -694
rect -527 -728 -493 -694
rect -459 -728 -425 -694
rect -391 -728 -357 -694
rect -323 -728 -289 -694
rect -255 -728 -221 -694
rect -187 -728 -153 -694
rect -119 -728 -85 -694
rect -51 -728 -17 -694
rect 17 -728 51 -694
rect 85 -728 119 -694
rect 153 -728 187 -694
rect 221 -728 255 -694
rect 289 -728 323 -694
rect 357 -728 391 -694
rect 425 -728 459 -694
rect 493 -728 527 -694
rect 561 -728 595 -694
rect 629 -728 663 -694
rect 697 -728 731 -694
rect 765 -728 799 -694
rect 833 -728 867 -694
rect 901 -728 935 -694
rect 969 -728 1003 -694
rect 1037 -728 1071 -694
rect 1105 -728 1139 -694
rect 1173 -728 1207 -694
rect 1241 -728 1275 -694
rect 1309 -728 1343 -694
rect 1377 -728 1411 -694
rect 1445 -728 1479 -694
rect 1513 -728 1547 -694
rect 1581 -728 1615 -694
rect 1649 -728 1683 -694
rect 1717 -728 1751 -694
rect 1785 -728 1819 -694
rect 1853 -728 1887 -694
rect 1921 -728 1955 -694
rect 1989 -728 2023 -694
rect 2057 -728 2091 -694
rect 2125 -728 2159 -694
rect 2193 -728 2227 -694
rect 2261 -728 2295 -694
rect 2329 -728 2363 -694
rect 2397 -728 2431 -694
rect 2465 -728 2499 -694
rect 2533 -728 2567 -694
rect 2601 -728 2635 -694
rect 2669 -728 2703 -694
rect 2737 -728 2771 -694
rect 2805 -728 2839 -694
rect 2873 -728 2907 -694
rect 2941 -728 2975 -694
rect 3009 -728 3043 -694
rect 3077 -728 3111 -694
rect 3145 -728 3179 -694
rect 3213 -728 3311 -694
<< viali >>
rect -3098 556 -3064 590
rect -2940 556 -2906 590
rect -2782 556 -2748 590
rect -2624 556 -2590 590
rect -2466 556 -2432 590
rect -2308 556 -2274 590
rect -2150 556 -2116 590
rect -1992 556 -1958 590
rect -1834 556 -1800 590
rect -1676 556 -1642 590
rect -1518 556 -1484 590
rect -1360 556 -1326 590
rect -1202 556 -1168 590
rect -1044 556 -1010 590
rect -886 556 -852 590
rect -728 556 -694 590
rect -570 556 -536 590
rect -412 556 -378 590
rect -254 556 -220 590
rect -96 556 -62 590
rect 62 556 96 590
rect 220 556 254 590
rect 378 556 412 590
rect 536 556 570 590
rect 694 556 728 590
rect 852 556 886 590
rect 1010 556 1044 590
rect 1168 556 1202 590
rect 1326 556 1360 590
rect 1484 556 1518 590
rect 1642 556 1676 590
rect 1800 556 1834 590
rect 1958 556 1992 590
rect 2116 556 2150 590
rect 2274 556 2308 590
rect 2432 556 2466 590
rect 2590 556 2624 590
rect 2748 556 2782 590
rect 2906 556 2940 590
rect 3064 556 3098 590
rect -3177 469 -3143 471
rect -3177 437 -3143 469
rect -3177 367 -3143 399
rect -3177 365 -3143 367
rect -3019 469 -2985 471
rect -3019 437 -2985 469
rect -3019 367 -2985 399
rect -3019 365 -2985 367
rect -2861 469 -2827 471
rect -2861 437 -2827 469
rect -2861 367 -2827 399
rect -2861 365 -2827 367
rect -2703 469 -2669 471
rect -2703 437 -2669 469
rect -2703 367 -2669 399
rect -2703 365 -2669 367
rect -2545 469 -2511 471
rect -2545 437 -2511 469
rect -2545 367 -2511 399
rect -2545 365 -2511 367
rect -2387 469 -2353 471
rect -2387 437 -2353 469
rect -2387 367 -2353 399
rect -2387 365 -2353 367
rect -2229 469 -2195 471
rect -2229 437 -2195 469
rect -2229 367 -2195 399
rect -2229 365 -2195 367
rect -2071 469 -2037 471
rect -2071 437 -2037 469
rect -2071 367 -2037 399
rect -2071 365 -2037 367
rect -1913 469 -1879 471
rect -1913 437 -1879 469
rect -1913 367 -1879 399
rect -1913 365 -1879 367
rect -1755 469 -1721 471
rect -1755 437 -1721 469
rect -1755 367 -1721 399
rect -1755 365 -1721 367
rect -1597 469 -1563 471
rect -1597 437 -1563 469
rect -1597 367 -1563 399
rect -1597 365 -1563 367
rect -1439 469 -1405 471
rect -1439 437 -1405 469
rect -1439 367 -1405 399
rect -1439 365 -1405 367
rect -1281 469 -1247 471
rect -1281 437 -1247 469
rect -1281 367 -1247 399
rect -1281 365 -1247 367
rect -1123 469 -1089 471
rect -1123 437 -1089 469
rect -1123 367 -1089 399
rect -1123 365 -1089 367
rect -965 469 -931 471
rect -965 437 -931 469
rect -965 367 -931 399
rect -965 365 -931 367
rect -807 469 -773 471
rect -807 437 -773 469
rect -807 367 -773 399
rect -807 365 -773 367
rect -649 469 -615 471
rect -649 437 -615 469
rect -649 367 -615 399
rect -649 365 -615 367
rect -491 469 -457 471
rect -491 437 -457 469
rect -491 367 -457 399
rect -491 365 -457 367
rect -333 469 -299 471
rect -333 437 -299 469
rect -333 367 -299 399
rect -333 365 -299 367
rect -175 469 -141 471
rect -175 437 -141 469
rect -175 367 -141 399
rect -175 365 -141 367
rect -17 469 17 471
rect -17 437 17 469
rect -17 367 17 399
rect -17 365 17 367
rect 141 469 175 471
rect 141 437 175 469
rect 141 367 175 399
rect 141 365 175 367
rect 299 469 333 471
rect 299 437 333 469
rect 299 367 333 399
rect 299 365 333 367
rect 457 469 491 471
rect 457 437 491 469
rect 457 367 491 399
rect 457 365 491 367
rect 615 469 649 471
rect 615 437 649 469
rect 615 367 649 399
rect 615 365 649 367
rect 773 469 807 471
rect 773 437 807 469
rect 773 367 807 399
rect 773 365 807 367
rect 931 469 965 471
rect 931 437 965 469
rect 931 367 965 399
rect 931 365 965 367
rect 1089 469 1123 471
rect 1089 437 1123 469
rect 1089 367 1123 399
rect 1089 365 1123 367
rect 1247 469 1281 471
rect 1247 437 1281 469
rect 1247 367 1281 399
rect 1247 365 1281 367
rect 1405 469 1439 471
rect 1405 437 1439 469
rect 1405 367 1439 399
rect 1405 365 1439 367
rect 1563 469 1597 471
rect 1563 437 1597 469
rect 1563 367 1597 399
rect 1563 365 1597 367
rect 1721 469 1755 471
rect 1721 437 1755 469
rect 1721 367 1755 399
rect 1721 365 1755 367
rect 1879 469 1913 471
rect 1879 437 1913 469
rect 1879 367 1913 399
rect 1879 365 1913 367
rect 2037 469 2071 471
rect 2037 437 2071 469
rect 2037 367 2071 399
rect 2037 365 2071 367
rect 2195 469 2229 471
rect 2195 437 2229 469
rect 2195 367 2229 399
rect 2195 365 2229 367
rect 2353 469 2387 471
rect 2353 437 2387 469
rect 2353 367 2387 399
rect 2353 365 2387 367
rect 2511 469 2545 471
rect 2511 437 2545 469
rect 2511 367 2545 399
rect 2511 365 2545 367
rect 2669 469 2703 471
rect 2669 437 2703 469
rect 2669 367 2703 399
rect 2669 365 2703 367
rect 2827 469 2861 471
rect 2827 437 2861 469
rect 2827 367 2861 399
rect 2827 365 2861 367
rect 2985 469 3019 471
rect 2985 437 3019 469
rect 2985 367 3019 399
rect 2985 365 3019 367
rect 3143 469 3177 471
rect 3143 437 3177 469
rect 3143 367 3177 399
rect 3143 365 3177 367
rect -3098 246 -3064 280
rect -2940 246 -2906 280
rect -2782 246 -2748 280
rect -2624 246 -2590 280
rect -2466 246 -2432 280
rect -2308 246 -2274 280
rect -2150 246 -2116 280
rect -1992 246 -1958 280
rect -1834 246 -1800 280
rect -1676 246 -1642 280
rect -1518 246 -1484 280
rect -1360 246 -1326 280
rect -1202 246 -1168 280
rect -1044 246 -1010 280
rect -886 246 -852 280
rect -728 246 -694 280
rect -570 246 -536 280
rect -412 246 -378 280
rect -254 246 -220 280
rect -96 246 -62 280
rect 62 246 96 280
rect 220 246 254 280
rect 378 246 412 280
rect 536 246 570 280
rect 694 246 728 280
rect 852 246 886 280
rect 1010 246 1044 280
rect 1168 246 1202 280
rect 1326 246 1360 280
rect 1484 246 1518 280
rect 1642 246 1676 280
rect 1800 246 1834 280
rect 1958 246 1992 280
rect 2116 246 2150 280
rect 2274 246 2308 280
rect 2432 246 2466 280
rect 2590 246 2624 280
rect 2748 246 2782 280
rect 2906 246 2940 280
rect 3064 246 3098 280
rect -3098 138 -3064 172
rect -2940 138 -2906 172
rect -2782 138 -2748 172
rect -2624 138 -2590 172
rect -2466 138 -2432 172
rect -2308 138 -2274 172
rect -2150 138 -2116 172
rect -1992 138 -1958 172
rect -1834 138 -1800 172
rect -1676 138 -1642 172
rect -1518 138 -1484 172
rect -1360 138 -1326 172
rect -1202 138 -1168 172
rect -1044 138 -1010 172
rect -886 138 -852 172
rect -728 138 -694 172
rect -570 138 -536 172
rect -412 138 -378 172
rect -254 138 -220 172
rect -96 138 -62 172
rect 62 138 96 172
rect 220 138 254 172
rect 378 138 412 172
rect 536 138 570 172
rect 694 138 728 172
rect 852 138 886 172
rect 1010 138 1044 172
rect 1168 138 1202 172
rect 1326 138 1360 172
rect 1484 138 1518 172
rect 1642 138 1676 172
rect 1800 138 1834 172
rect 1958 138 1992 172
rect 2116 138 2150 172
rect 2274 138 2308 172
rect 2432 138 2466 172
rect 2590 138 2624 172
rect 2748 138 2782 172
rect 2906 138 2940 172
rect 3064 138 3098 172
rect -3177 51 -3143 53
rect -3177 19 -3143 51
rect -3177 -51 -3143 -19
rect -3177 -53 -3143 -51
rect -3019 51 -2985 53
rect -3019 19 -2985 51
rect -3019 -51 -2985 -19
rect -3019 -53 -2985 -51
rect -2861 51 -2827 53
rect -2861 19 -2827 51
rect -2861 -51 -2827 -19
rect -2861 -53 -2827 -51
rect -2703 51 -2669 53
rect -2703 19 -2669 51
rect -2703 -51 -2669 -19
rect -2703 -53 -2669 -51
rect -2545 51 -2511 53
rect -2545 19 -2511 51
rect -2545 -51 -2511 -19
rect -2545 -53 -2511 -51
rect -2387 51 -2353 53
rect -2387 19 -2353 51
rect -2387 -51 -2353 -19
rect -2387 -53 -2353 -51
rect -2229 51 -2195 53
rect -2229 19 -2195 51
rect -2229 -51 -2195 -19
rect -2229 -53 -2195 -51
rect -2071 51 -2037 53
rect -2071 19 -2037 51
rect -2071 -51 -2037 -19
rect -2071 -53 -2037 -51
rect -1913 51 -1879 53
rect -1913 19 -1879 51
rect -1913 -51 -1879 -19
rect -1913 -53 -1879 -51
rect -1755 51 -1721 53
rect -1755 19 -1721 51
rect -1755 -51 -1721 -19
rect -1755 -53 -1721 -51
rect -1597 51 -1563 53
rect -1597 19 -1563 51
rect -1597 -51 -1563 -19
rect -1597 -53 -1563 -51
rect -1439 51 -1405 53
rect -1439 19 -1405 51
rect -1439 -51 -1405 -19
rect -1439 -53 -1405 -51
rect -1281 51 -1247 53
rect -1281 19 -1247 51
rect -1281 -51 -1247 -19
rect -1281 -53 -1247 -51
rect -1123 51 -1089 53
rect -1123 19 -1089 51
rect -1123 -51 -1089 -19
rect -1123 -53 -1089 -51
rect -965 51 -931 53
rect -965 19 -931 51
rect -965 -51 -931 -19
rect -965 -53 -931 -51
rect -807 51 -773 53
rect -807 19 -773 51
rect -807 -51 -773 -19
rect -807 -53 -773 -51
rect -649 51 -615 53
rect -649 19 -615 51
rect -649 -51 -615 -19
rect -649 -53 -615 -51
rect -491 51 -457 53
rect -491 19 -457 51
rect -491 -51 -457 -19
rect -491 -53 -457 -51
rect -333 51 -299 53
rect -333 19 -299 51
rect -333 -51 -299 -19
rect -333 -53 -299 -51
rect -175 51 -141 53
rect -175 19 -141 51
rect -175 -51 -141 -19
rect -175 -53 -141 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 141 51 175 53
rect 141 19 175 51
rect 141 -51 175 -19
rect 141 -53 175 -51
rect 299 51 333 53
rect 299 19 333 51
rect 299 -51 333 -19
rect 299 -53 333 -51
rect 457 51 491 53
rect 457 19 491 51
rect 457 -51 491 -19
rect 457 -53 491 -51
rect 615 51 649 53
rect 615 19 649 51
rect 615 -51 649 -19
rect 615 -53 649 -51
rect 773 51 807 53
rect 773 19 807 51
rect 773 -51 807 -19
rect 773 -53 807 -51
rect 931 51 965 53
rect 931 19 965 51
rect 931 -51 965 -19
rect 931 -53 965 -51
rect 1089 51 1123 53
rect 1089 19 1123 51
rect 1089 -51 1123 -19
rect 1089 -53 1123 -51
rect 1247 51 1281 53
rect 1247 19 1281 51
rect 1247 -51 1281 -19
rect 1247 -53 1281 -51
rect 1405 51 1439 53
rect 1405 19 1439 51
rect 1405 -51 1439 -19
rect 1405 -53 1439 -51
rect 1563 51 1597 53
rect 1563 19 1597 51
rect 1563 -51 1597 -19
rect 1563 -53 1597 -51
rect 1721 51 1755 53
rect 1721 19 1755 51
rect 1721 -51 1755 -19
rect 1721 -53 1755 -51
rect 1879 51 1913 53
rect 1879 19 1913 51
rect 1879 -51 1913 -19
rect 1879 -53 1913 -51
rect 2037 51 2071 53
rect 2037 19 2071 51
rect 2037 -51 2071 -19
rect 2037 -53 2071 -51
rect 2195 51 2229 53
rect 2195 19 2229 51
rect 2195 -51 2229 -19
rect 2195 -53 2229 -51
rect 2353 51 2387 53
rect 2353 19 2387 51
rect 2353 -51 2387 -19
rect 2353 -53 2387 -51
rect 2511 51 2545 53
rect 2511 19 2545 51
rect 2511 -51 2545 -19
rect 2511 -53 2545 -51
rect 2669 51 2703 53
rect 2669 19 2703 51
rect 2669 -51 2703 -19
rect 2669 -53 2703 -51
rect 2827 51 2861 53
rect 2827 19 2861 51
rect 2827 -51 2861 -19
rect 2827 -53 2861 -51
rect 2985 51 3019 53
rect 2985 19 3019 51
rect 2985 -51 3019 -19
rect 2985 -53 3019 -51
rect 3143 51 3177 53
rect 3143 19 3177 51
rect 3143 -51 3177 -19
rect 3143 -53 3177 -51
rect -3098 -172 -3064 -138
rect -2940 -172 -2906 -138
rect -2782 -172 -2748 -138
rect -2624 -172 -2590 -138
rect -2466 -172 -2432 -138
rect -2308 -172 -2274 -138
rect -2150 -172 -2116 -138
rect -1992 -172 -1958 -138
rect -1834 -172 -1800 -138
rect -1676 -172 -1642 -138
rect -1518 -172 -1484 -138
rect -1360 -172 -1326 -138
rect -1202 -172 -1168 -138
rect -1044 -172 -1010 -138
rect -886 -172 -852 -138
rect -728 -172 -694 -138
rect -570 -172 -536 -138
rect -412 -172 -378 -138
rect -254 -172 -220 -138
rect -96 -172 -62 -138
rect 62 -172 96 -138
rect 220 -172 254 -138
rect 378 -172 412 -138
rect 536 -172 570 -138
rect 694 -172 728 -138
rect 852 -172 886 -138
rect 1010 -172 1044 -138
rect 1168 -172 1202 -138
rect 1326 -172 1360 -138
rect 1484 -172 1518 -138
rect 1642 -172 1676 -138
rect 1800 -172 1834 -138
rect 1958 -172 1992 -138
rect 2116 -172 2150 -138
rect 2274 -172 2308 -138
rect 2432 -172 2466 -138
rect 2590 -172 2624 -138
rect 2748 -172 2782 -138
rect 2906 -172 2940 -138
rect 3064 -172 3098 -138
rect -3098 -280 -3064 -246
rect -2940 -280 -2906 -246
rect -2782 -280 -2748 -246
rect -2624 -280 -2590 -246
rect -2466 -280 -2432 -246
rect -2308 -280 -2274 -246
rect -2150 -280 -2116 -246
rect -1992 -280 -1958 -246
rect -1834 -280 -1800 -246
rect -1676 -280 -1642 -246
rect -1518 -280 -1484 -246
rect -1360 -280 -1326 -246
rect -1202 -280 -1168 -246
rect -1044 -280 -1010 -246
rect -886 -280 -852 -246
rect -728 -280 -694 -246
rect -570 -280 -536 -246
rect -412 -280 -378 -246
rect -254 -280 -220 -246
rect -96 -280 -62 -246
rect 62 -280 96 -246
rect 220 -280 254 -246
rect 378 -280 412 -246
rect 536 -280 570 -246
rect 694 -280 728 -246
rect 852 -280 886 -246
rect 1010 -280 1044 -246
rect 1168 -280 1202 -246
rect 1326 -280 1360 -246
rect 1484 -280 1518 -246
rect 1642 -280 1676 -246
rect 1800 -280 1834 -246
rect 1958 -280 1992 -246
rect 2116 -280 2150 -246
rect 2274 -280 2308 -246
rect 2432 -280 2466 -246
rect 2590 -280 2624 -246
rect 2748 -280 2782 -246
rect 2906 -280 2940 -246
rect 3064 -280 3098 -246
rect -3177 -367 -3143 -365
rect -3177 -399 -3143 -367
rect -3177 -469 -3143 -437
rect -3177 -471 -3143 -469
rect -3019 -367 -2985 -365
rect -3019 -399 -2985 -367
rect -3019 -469 -2985 -437
rect -3019 -471 -2985 -469
rect -2861 -367 -2827 -365
rect -2861 -399 -2827 -367
rect -2861 -469 -2827 -437
rect -2861 -471 -2827 -469
rect -2703 -367 -2669 -365
rect -2703 -399 -2669 -367
rect -2703 -469 -2669 -437
rect -2703 -471 -2669 -469
rect -2545 -367 -2511 -365
rect -2545 -399 -2511 -367
rect -2545 -469 -2511 -437
rect -2545 -471 -2511 -469
rect -2387 -367 -2353 -365
rect -2387 -399 -2353 -367
rect -2387 -469 -2353 -437
rect -2387 -471 -2353 -469
rect -2229 -367 -2195 -365
rect -2229 -399 -2195 -367
rect -2229 -469 -2195 -437
rect -2229 -471 -2195 -469
rect -2071 -367 -2037 -365
rect -2071 -399 -2037 -367
rect -2071 -469 -2037 -437
rect -2071 -471 -2037 -469
rect -1913 -367 -1879 -365
rect -1913 -399 -1879 -367
rect -1913 -469 -1879 -437
rect -1913 -471 -1879 -469
rect -1755 -367 -1721 -365
rect -1755 -399 -1721 -367
rect -1755 -469 -1721 -437
rect -1755 -471 -1721 -469
rect -1597 -367 -1563 -365
rect -1597 -399 -1563 -367
rect -1597 -469 -1563 -437
rect -1597 -471 -1563 -469
rect -1439 -367 -1405 -365
rect -1439 -399 -1405 -367
rect -1439 -469 -1405 -437
rect -1439 -471 -1405 -469
rect -1281 -367 -1247 -365
rect -1281 -399 -1247 -367
rect -1281 -469 -1247 -437
rect -1281 -471 -1247 -469
rect -1123 -367 -1089 -365
rect -1123 -399 -1089 -367
rect -1123 -469 -1089 -437
rect -1123 -471 -1089 -469
rect -965 -367 -931 -365
rect -965 -399 -931 -367
rect -965 -469 -931 -437
rect -965 -471 -931 -469
rect -807 -367 -773 -365
rect -807 -399 -773 -367
rect -807 -469 -773 -437
rect -807 -471 -773 -469
rect -649 -367 -615 -365
rect -649 -399 -615 -367
rect -649 -469 -615 -437
rect -649 -471 -615 -469
rect -491 -367 -457 -365
rect -491 -399 -457 -367
rect -491 -469 -457 -437
rect -491 -471 -457 -469
rect -333 -367 -299 -365
rect -333 -399 -299 -367
rect -333 -469 -299 -437
rect -333 -471 -299 -469
rect -175 -367 -141 -365
rect -175 -399 -141 -367
rect -175 -469 -141 -437
rect -175 -471 -141 -469
rect -17 -367 17 -365
rect -17 -399 17 -367
rect -17 -469 17 -437
rect -17 -471 17 -469
rect 141 -367 175 -365
rect 141 -399 175 -367
rect 141 -469 175 -437
rect 141 -471 175 -469
rect 299 -367 333 -365
rect 299 -399 333 -367
rect 299 -469 333 -437
rect 299 -471 333 -469
rect 457 -367 491 -365
rect 457 -399 491 -367
rect 457 -469 491 -437
rect 457 -471 491 -469
rect 615 -367 649 -365
rect 615 -399 649 -367
rect 615 -469 649 -437
rect 615 -471 649 -469
rect 773 -367 807 -365
rect 773 -399 807 -367
rect 773 -469 807 -437
rect 773 -471 807 -469
rect 931 -367 965 -365
rect 931 -399 965 -367
rect 931 -469 965 -437
rect 931 -471 965 -469
rect 1089 -367 1123 -365
rect 1089 -399 1123 -367
rect 1089 -469 1123 -437
rect 1089 -471 1123 -469
rect 1247 -367 1281 -365
rect 1247 -399 1281 -367
rect 1247 -469 1281 -437
rect 1247 -471 1281 -469
rect 1405 -367 1439 -365
rect 1405 -399 1439 -367
rect 1405 -469 1439 -437
rect 1405 -471 1439 -469
rect 1563 -367 1597 -365
rect 1563 -399 1597 -367
rect 1563 -469 1597 -437
rect 1563 -471 1597 -469
rect 1721 -367 1755 -365
rect 1721 -399 1755 -367
rect 1721 -469 1755 -437
rect 1721 -471 1755 -469
rect 1879 -367 1913 -365
rect 1879 -399 1913 -367
rect 1879 -469 1913 -437
rect 1879 -471 1913 -469
rect 2037 -367 2071 -365
rect 2037 -399 2071 -367
rect 2037 -469 2071 -437
rect 2037 -471 2071 -469
rect 2195 -367 2229 -365
rect 2195 -399 2229 -367
rect 2195 -469 2229 -437
rect 2195 -471 2229 -469
rect 2353 -367 2387 -365
rect 2353 -399 2387 -367
rect 2353 -469 2387 -437
rect 2353 -471 2387 -469
rect 2511 -367 2545 -365
rect 2511 -399 2545 -367
rect 2511 -469 2545 -437
rect 2511 -471 2545 -469
rect 2669 -367 2703 -365
rect 2669 -399 2703 -367
rect 2669 -469 2703 -437
rect 2669 -471 2703 -469
rect 2827 -367 2861 -365
rect 2827 -399 2861 -367
rect 2827 -469 2861 -437
rect 2827 -471 2861 -469
rect 2985 -367 3019 -365
rect 2985 -399 3019 -367
rect 2985 -469 3019 -437
rect 2985 -471 3019 -469
rect 3143 -367 3177 -365
rect 3143 -399 3177 -367
rect 3143 -469 3177 -437
rect 3143 -471 3177 -469
rect -3098 -590 -3064 -556
rect -2940 -590 -2906 -556
rect -2782 -590 -2748 -556
rect -2624 -590 -2590 -556
rect -2466 -590 -2432 -556
rect -2308 -590 -2274 -556
rect -2150 -590 -2116 -556
rect -1992 -590 -1958 -556
rect -1834 -590 -1800 -556
rect -1676 -590 -1642 -556
rect -1518 -590 -1484 -556
rect -1360 -590 -1326 -556
rect -1202 -590 -1168 -556
rect -1044 -590 -1010 -556
rect -886 -590 -852 -556
rect -728 -590 -694 -556
rect -570 -590 -536 -556
rect -412 -590 -378 -556
rect -254 -590 -220 -556
rect -96 -590 -62 -556
rect 62 -590 96 -556
rect 220 -590 254 -556
rect 378 -590 412 -556
rect 536 -590 570 -556
rect 694 -590 728 -556
rect 852 -590 886 -556
rect 1010 -590 1044 -556
rect 1168 -590 1202 -556
rect 1326 -590 1360 -556
rect 1484 -590 1518 -556
rect 1642 -590 1676 -556
rect 1800 -590 1834 -556
rect 1958 -590 1992 -556
rect 2116 -590 2150 -556
rect 2274 -590 2308 -556
rect 2432 -590 2466 -556
rect 2590 -590 2624 -556
rect 2748 -590 2782 -556
rect 2906 -590 2940 -556
rect 3064 -590 3098 -556
<< metal1 >>
rect -3127 590 -3035 596
rect -3127 556 -3098 590
rect -3064 556 -3035 590
rect -3127 550 -3035 556
rect -2969 590 -2877 596
rect -2969 556 -2940 590
rect -2906 556 -2877 590
rect -2969 550 -2877 556
rect -2811 590 -2719 596
rect -2811 556 -2782 590
rect -2748 556 -2719 590
rect -2811 550 -2719 556
rect -2653 590 -2561 596
rect -2653 556 -2624 590
rect -2590 556 -2561 590
rect -2653 550 -2561 556
rect -2495 590 -2403 596
rect -2495 556 -2466 590
rect -2432 556 -2403 590
rect -2495 550 -2403 556
rect -2337 590 -2245 596
rect -2337 556 -2308 590
rect -2274 556 -2245 590
rect -2337 550 -2245 556
rect -2179 590 -2087 596
rect -2179 556 -2150 590
rect -2116 556 -2087 590
rect -2179 550 -2087 556
rect -2021 590 -1929 596
rect -2021 556 -1992 590
rect -1958 556 -1929 590
rect -2021 550 -1929 556
rect -1863 590 -1771 596
rect -1863 556 -1834 590
rect -1800 556 -1771 590
rect -1863 550 -1771 556
rect -1705 590 -1613 596
rect -1705 556 -1676 590
rect -1642 556 -1613 590
rect -1705 550 -1613 556
rect -1547 590 -1455 596
rect -1547 556 -1518 590
rect -1484 556 -1455 590
rect -1547 550 -1455 556
rect -1389 590 -1297 596
rect -1389 556 -1360 590
rect -1326 556 -1297 590
rect -1389 550 -1297 556
rect -1231 590 -1139 596
rect -1231 556 -1202 590
rect -1168 556 -1139 590
rect -1231 550 -1139 556
rect -1073 590 -981 596
rect -1073 556 -1044 590
rect -1010 556 -981 590
rect -1073 550 -981 556
rect -915 590 -823 596
rect -915 556 -886 590
rect -852 556 -823 590
rect -915 550 -823 556
rect -757 590 -665 596
rect -757 556 -728 590
rect -694 556 -665 590
rect -757 550 -665 556
rect -599 590 -507 596
rect -599 556 -570 590
rect -536 556 -507 590
rect -599 550 -507 556
rect -441 590 -349 596
rect -441 556 -412 590
rect -378 556 -349 590
rect -441 550 -349 556
rect -283 590 -191 596
rect -283 556 -254 590
rect -220 556 -191 590
rect -283 550 -191 556
rect -125 590 -33 596
rect -125 556 -96 590
rect -62 556 -33 590
rect -125 550 -33 556
rect 33 590 125 596
rect 33 556 62 590
rect 96 556 125 590
rect 33 550 125 556
rect 191 590 283 596
rect 191 556 220 590
rect 254 556 283 590
rect 191 550 283 556
rect 349 590 441 596
rect 349 556 378 590
rect 412 556 441 590
rect 349 550 441 556
rect 507 590 599 596
rect 507 556 536 590
rect 570 556 599 590
rect 507 550 599 556
rect 665 590 757 596
rect 665 556 694 590
rect 728 556 757 590
rect 665 550 757 556
rect 823 590 915 596
rect 823 556 852 590
rect 886 556 915 590
rect 823 550 915 556
rect 981 590 1073 596
rect 981 556 1010 590
rect 1044 556 1073 590
rect 981 550 1073 556
rect 1139 590 1231 596
rect 1139 556 1168 590
rect 1202 556 1231 590
rect 1139 550 1231 556
rect 1297 590 1389 596
rect 1297 556 1326 590
rect 1360 556 1389 590
rect 1297 550 1389 556
rect 1455 590 1547 596
rect 1455 556 1484 590
rect 1518 556 1547 590
rect 1455 550 1547 556
rect 1613 590 1705 596
rect 1613 556 1642 590
rect 1676 556 1705 590
rect 1613 550 1705 556
rect 1771 590 1863 596
rect 1771 556 1800 590
rect 1834 556 1863 590
rect 1771 550 1863 556
rect 1929 590 2021 596
rect 1929 556 1958 590
rect 1992 556 2021 590
rect 1929 550 2021 556
rect 2087 590 2179 596
rect 2087 556 2116 590
rect 2150 556 2179 590
rect 2087 550 2179 556
rect 2245 590 2337 596
rect 2245 556 2274 590
rect 2308 556 2337 590
rect 2245 550 2337 556
rect 2403 590 2495 596
rect 2403 556 2432 590
rect 2466 556 2495 590
rect 2403 550 2495 556
rect 2561 590 2653 596
rect 2561 556 2590 590
rect 2624 556 2653 590
rect 2561 550 2653 556
rect 2719 590 2811 596
rect 2719 556 2748 590
rect 2782 556 2811 590
rect 2719 550 2811 556
rect 2877 590 2969 596
rect 2877 556 2906 590
rect 2940 556 2969 590
rect 2877 550 2969 556
rect 3035 590 3127 596
rect 3035 556 3064 590
rect 3098 556 3127 590
rect 3035 550 3127 556
rect -3183 471 -3137 518
rect -3183 437 -3177 471
rect -3143 437 -3137 471
rect -3183 399 -3137 437
rect -3183 365 -3177 399
rect -3143 365 -3137 399
rect -3183 318 -3137 365
rect -3025 471 -2979 518
rect -3025 437 -3019 471
rect -2985 437 -2979 471
rect -3025 399 -2979 437
rect -3025 365 -3019 399
rect -2985 365 -2979 399
rect -3025 318 -2979 365
rect -2867 471 -2821 518
rect -2867 437 -2861 471
rect -2827 437 -2821 471
rect -2867 399 -2821 437
rect -2867 365 -2861 399
rect -2827 365 -2821 399
rect -2867 318 -2821 365
rect -2709 471 -2663 518
rect -2709 437 -2703 471
rect -2669 437 -2663 471
rect -2709 399 -2663 437
rect -2709 365 -2703 399
rect -2669 365 -2663 399
rect -2709 318 -2663 365
rect -2551 471 -2505 518
rect -2551 437 -2545 471
rect -2511 437 -2505 471
rect -2551 399 -2505 437
rect -2551 365 -2545 399
rect -2511 365 -2505 399
rect -2551 318 -2505 365
rect -2393 471 -2347 518
rect -2393 437 -2387 471
rect -2353 437 -2347 471
rect -2393 399 -2347 437
rect -2393 365 -2387 399
rect -2353 365 -2347 399
rect -2393 318 -2347 365
rect -2235 471 -2189 518
rect -2235 437 -2229 471
rect -2195 437 -2189 471
rect -2235 399 -2189 437
rect -2235 365 -2229 399
rect -2195 365 -2189 399
rect -2235 318 -2189 365
rect -2077 471 -2031 518
rect -2077 437 -2071 471
rect -2037 437 -2031 471
rect -2077 399 -2031 437
rect -2077 365 -2071 399
rect -2037 365 -2031 399
rect -2077 318 -2031 365
rect -1919 471 -1873 518
rect -1919 437 -1913 471
rect -1879 437 -1873 471
rect -1919 399 -1873 437
rect -1919 365 -1913 399
rect -1879 365 -1873 399
rect -1919 318 -1873 365
rect -1761 471 -1715 518
rect -1761 437 -1755 471
rect -1721 437 -1715 471
rect -1761 399 -1715 437
rect -1761 365 -1755 399
rect -1721 365 -1715 399
rect -1761 318 -1715 365
rect -1603 471 -1557 518
rect -1603 437 -1597 471
rect -1563 437 -1557 471
rect -1603 399 -1557 437
rect -1603 365 -1597 399
rect -1563 365 -1557 399
rect -1603 318 -1557 365
rect -1445 471 -1399 518
rect -1445 437 -1439 471
rect -1405 437 -1399 471
rect -1445 399 -1399 437
rect -1445 365 -1439 399
rect -1405 365 -1399 399
rect -1445 318 -1399 365
rect -1287 471 -1241 518
rect -1287 437 -1281 471
rect -1247 437 -1241 471
rect -1287 399 -1241 437
rect -1287 365 -1281 399
rect -1247 365 -1241 399
rect -1287 318 -1241 365
rect -1129 471 -1083 518
rect -1129 437 -1123 471
rect -1089 437 -1083 471
rect -1129 399 -1083 437
rect -1129 365 -1123 399
rect -1089 365 -1083 399
rect -1129 318 -1083 365
rect -971 471 -925 518
rect -971 437 -965 471
rect -931 437 -925 471
rect -971 399 -925 437
rect -971 365 -965 399
rect -931 365 -925 399
rect -971 318 -925 365
rect -813 471 -767 518
rect -813 437 -807 471
rect -773 437 -767 471
rect -813 399 -767 437
rect -813 365 -807 399
rect -773 365 -767 399
rect -813 318 -767 365
rect -655 471 -609 518
rect -655 437 -649 471
rect -615 437 -609 471
rect -655 399 -609 437
rect -655 365 -649 399
rect -615 365 -609 399
rect -655 318 -609 365
rect -497 471 -451 518
rect -497 437 -491 471
rect -457 437 -451 471
rect -497 399 -451 437
rect -497 365 -491 399
rect -457 365 -451 399
rect -497 318 -451 365
rect -339 471 -293 518
rect -339 437 -333 471
rect -299 437 -293 471
rect -339 399 -293 437
rect -339 365 -333 399
rect -299 365 -293 399
rect -339 318 -293 365
rect -181 471 -135 518
rect -181 437 -175 471
rect -141 437 -135 471
rect -181 399 -135 437
rect -181 365 -175 399
rect -141 365 -135 399
rect -181 318 -135 365
rect -23 471 23 518
rect -23 437 -17 471
rect 17 437 23 471
rect -23 399 23 437
rect -23 365 -17 399
rect 17 365 23 399
rect -23 318 23 365
rect 135 471 181 518
rect 135 437 141 471
rect 175 437 181 471
rect 135 399 181 437
rect 135 365 141 399
rect 175 365 181 399
rect 135 318 181 365
rect 293 471 339 518
rect 293 437 299 471
rect 333 437 339 471
rect 293 399 339 437
rect 293 365 299 399
rect 333 365 339 399
rect 293 318 339 365
rect 451 471 497 518
rect 451 437 457 471
rect 491 437 497 471
rect 451 399 497 437
rect 451 365 457 399
rect 491 365 497 399
rect 451 318 497 365
rect 609 471 655 518
rect 609 437 615 471
rect 649 437 655 471
rect 609 399 655 437
rect 609 365 615 399
rect 649 365 655 399
rect 609 318 655 365
rect 767 471 813 518
rect 767 437 773 471
rect 807 437 813 471
rect 767 399 813 437
rect 767 365 773 399
rect 807 365 813 399
rect 767 318 813 365
rect 925 471 971 518
rect 925 437 931 471
rect 965 437 971 471
rect 925 399 971 437
rect 925 365 931 399
rect 965 365 971 399
rect 925 318 971 365
rect 1083 471 1129 518
rect 1083 437 1089 471
rect 1123 437 1129 471
rect 1083 399 1129 437
rect 1083 365 1089 399
rect 1123 365 1129 399
rect 1083 318 1129 365
rect 1241 471 1287 518
rect 1241 437 1247 471
rect 1281 437 1287 471
rect 1241 399 1287 437
rect 1241 365 1247 399
rect 1281 365 1287 399
rect 1241 318 1287 365
rect 1399 471 1445 518
rect 1399 437 1405 471
rect 1439 437 1445 471
rect 1399 399 1445 437
rect 1399 365 1405 399
rect 1439 365 1445 399
rect 1399 318 1445 365
rect 1557 471 1603 518
rect 1557 437 1563 471
rect 1597 437 1603 471
rect 1557 399 1603 437
rect 1557 365 1563 399
rect 1597 365 1603 399
rect 1557 318 1603 365
rect 1715 471 1761 518
rect 1715 437 1721 471
rect 1755 437 1761 471
rect 1715 399 1761 437
rect 1715 365 1721 399
rect 1755 365 1761 399
rect 1715 318 1761 365
rect 1873 471 1919 518
rect 1873 437 1879 471
rect 1913 437 1919 471
rect 1873 399 1919 437
rect 1873 365 1879 399
rect 1913 365 1919 399
rect 1873 318 1919 365
rect 2031 471 2077 518
rect 2031 437 2037 471
rect 2071 437 2077 471
rect 2031 399 2077 437
rect 2031 365 2037 399
rect 2071 365 2077 399
rect 2031 318 2077 365
rect 2189 471 2235 518
rect 2189 437 2195 471
rect 2229 437 2235 471
rect 2189 399 2235 437
rect 2189 365 2195 399
rect 2229 365 2235 399
rect 2189 318 2235 365
rect 2347 471 2393 518
rect 2347 437 2353 471
rect 2387 437 2393 471
rect 2347 399 2393 437
rect 2347 365 2353 399
rect 2387 365 2393 399
rect 2347 318 2393 365
rect 2505 471 2551 518
rect 2505 437 2511 471
rect 2545 437 2551 471
rect 2505 399 2551 437
rect 2505 365 2511 399
rect 2545 365 2551 399
rect 2505 318 2551 365
rect 2663 471 2709 518
rect 2663 437 2669 471
rect 2703 437 2709 471
rect 2663 399 2709 437
rect 2663 365 2669 399
rect 2703 365 2709 399
rect 2663 318 2709 365
rect 2821 471 2867 518
rect 2821 437 2827 471
rect 2861 437 2867 471
rect 2821 399 2867 437
rect 2821 365 2827 399
rect 2861 365 2867 399
rect 2821 318 2867 365
rect 2979 471 3025 518
rect 2979 437 2985 471
rect 3019 437 3025 471
rect 2979 399 3025 437
rect 2979 365 2985 399
rect 3019 365 3025 399
rect 2979 318 3025 365
rect 3137 471 3183 518
rect 3137 437 3143 471
rect 3177 437 3183 471
rect 3137 399 3183 437
rect 3137 365 3143 399
rect 3177 365 3183 399
rect 3137 318 3183 365
rect -3127 280 -3035 286
rect -3127 246 -3098 280
rect -3064 246 -3035 280
rect -3127 240 -3035 246
rect -2969 280 -2877 286
rect -2969 246 -2940 280
rect -2906 246 -2877 280
rect -2969 240 -2877 246
rect -2811 280 -2719 286
rect -2811 246 -2782 280
rect -2748 246 -2719 280
rect -2811 240 -2719 246
rect -2653 280 -2561 286
rect -2653 246 -2624 280
rect -2590 246 -2561 280
rect -2653 240 -2561 246
rect -2495 280 -2403 286
rect -2495 246 -2466 280
rect -2432 246 -2403 280
rect -2495 240 -2403 246
rect -2337 280 -2245 286
rect -2337 246 -2308 280
rect -2274 246 -2245 280
rect -2337 240 -2245 246
rect -2179 280 -2087 286
rect -2179 246 -2150 280
rect -2116 246 -2087 280
rect -2179 240 -2087 246
rect -2021 280 -1929 286
rect -2021 246 -1992 280
rect -1958 246 -1929 280
rect -2021 240 -1929 246
rect -1863 280 -1771 286
rect -1863 246 -1834 280
rect -1800 246 -1771 280
rect -1863 240 -1771 246
rect -1705 280 -1613 286
rect -1705 246 -1676 280
rect -1642 246 -1613 280
rect -1705 240 -1613 246
rect -1547 280 -1455 286
rect -1547 246 -1518 280
rect -1484 246 -1455 280
rect -1547 240 -1455 246
rect -1389 280 -1297 286
rect -1389 246 -1360 280
rect -1326 246 -1297 280
rect -1389 240 -1297 246
rect -1231 280 -1139 286
rect -1231 246 -1202 280
rect -1168 246 -1139 280
rect -1231 240 -1139 246
rect -1073 280 -981 286
rect -1073 246 -1044 280
rect -1010 246 -981 280
rect -1073 240 -981 246
rect -915 280 -823 286
rect -915 246 -886 280
rect -852 246 -823 280
rect -915 240 -823 246
rect -757 280 -665 286
rect -757 246 -728 280
rect -694 246 -665 280
rect -757 240 -665 246
rect -599 280 -507 286
rect -599 246 -570 280
rect -536 246 -507 280
rect -599 240 -507 246
rect -441 280 -349 286
rect -441 246 -412 280
rect -378 246 -349 280
rect -441 240 -349 246
rect -283 280 -191 286
rect -283 246 -254 280
rect -220 246 -191 280
rect -283 240 -191 246
rect -125 280 -33 286
rect -125 246 -96 280
rect -62 246 -33 280
rect -125 240 -33 246
rect 33 280 125 286
rect 33 246 62 280
rect 96 246 125 280
rect 33 240 125 246
rect 191 280 283 286
rect 191 246 220 280
rect 254 246 283 280
rect 191 240 283 246
rect 349 280 441 286
rect 349 246 378 280
rect 412 246 441 280
rect 349 240 441 246
rect 507 280 599 286
rect 507 246 536 280
rect 570 246 599 280
rect 507 240 599 246
rect 665 280 757 286
rect 665 246 694 280
rect 728 246 757 280
rect 665 240 757 246
rect 823 280 915 286
rect 823 246 852 280
rect 886 246 915 280
rect 823 240 915 246
rect 981 280 1073 286
rect 981 246 1010 280
rect 1044 246 1073 280
rect 981 240 1073 246
rect 1139 280 1231 286
rect 1139 246 1168 280
rect 1202 246 1231 280
rect 1139 240 1231 246
rect 1297 280 1389 286
rect 1297 246 1326 280
rect 1360 246 1389 280
rect 1297 240 1389 246
rect 1455 280 1547 286
rect 1455 246 1484 280
rect 1518 246 1547 280
rect 1455 240 1547 246
rect 1613 280 1705 286
rect 1613 246 1642 280
rect 1676 246 1705 280
rect 1613 240 1705 246
rect 1771 280 1863 286
rect 1771 246 1800 280
rect 1834 246 1863 280
rect 1771 240 1863 246
rect 1929 280 2021 286
rect 1929 246 1958 280
rect 1992 246 2021 280
rect 1929 240 2021 246
rect 2087 280 2179 286
rect 2087 246 2116 280
rect 2150 246 2179 280
rect 2087 240 2179 246
rect 2245 280 2337 286
rect 2245 246 2274 280
rect 2308 246 2337 280
rect 2245 240 2337 246
rect 2403 280 2495 286
rect 2403 246 2432 280
rect 2466 246 2495 280
rect 2403 240 2495 246
rect 2561 280 2653 286
rect 2561 246 2590 280
rect 2624 246 2653 280
rect 2561 240 2653 246
rect 2719 280 2811 286
rect 2719 246 2748 280
rect 2782 246 2811 280
rect 2719 240 2811 246
rect 2877 280 2969 286
rect 2877 246 2906 280
rect 2940 246 2969 280
rect 2877 240 2969 246
rect 3035 280 3127 286
rect 3035 246 3064 280
rect 3098 246 3127 280
rect 3035 240 3127 246
rect -3127 172 -3035 178
rect -3127 138 -3098 172
rect -3064 138 -3035 172
rect -3127 132 -3035 138
rect -2969 172 -2877 178
rect -2969 138 -2940 172
rect -2906 138 -2877 172
rect -2969 132 -2877 138
rect -2811 172 -2719 178
rect -2811 138 -2782 172
rect -2748 138 -2719 172
rect -2811 132 -2719 138
rect -2653 172 -2561 178
rect -2653 138 -2624 172
rect -2590 138 -2561 172
rect -2653 132 -2561 138
rect -2495 172 -2403 178
rect -2495 138 -2466 172
rect -2432 138 -2403 172
rect -2495 132 -2403 138
rect -2337 172 -2245 178
rect -2337 138 -2308 172
rect -2274 138 -2245 172
rect -2337 132 -2245 138
rect -2179 172 -2087 178
rect -2179 138 -2150 172
rect -2116 138 -2087 172
rect -2179 132 -2087 138
rect -2021 172 -1929 178
rect -2021 138 -1992 172
rect -1958 138 -1929 172
rect -2021 132 -1929 138
rect -1863 172 -1771 178
rect -1863 138 -1834 172
rect -1800 138 -1771 172
rect -1863 132 -1771 138
rect -1705 172 -1613 178
rect -1705 138 -1676 172
rect -1642 138 -1613 172
rect -1705 132 -1613 138
rect -1547 172 -1455 178
rect -1547 138 -1518 172
rect -1484 138 -1455 172
rect -1547 132 -1455 138
rect -1389 172 -1297 178
rect -1389 138 -1360 172
rect -1326 138 -1297 172
rect -1389 132 -1297 138
rect -1231 172 -1139 178
rect -1231 138 -1202 172
rect -1168 138 -1139 172
rect -1231 132 -1139 138
rect -1073 172 -981 178
rect -1073 138 -1044 172
rect -1010 138 -981 172
rect -1073 132 -981 138
rect -915 172 -823 178
rect -915 138 -886 172
rect -852 138 -823 172
rect -915 132 -823 138
rect -757 172 -665 178
rect -757 138 -728 172
rect -694 138 -665 172
rect -757 132 -665 138
rect -599 172 -507 178
rect -599 138 -570 172
rect -536 138 -507 172
rect -599 132 -507 138
rect -441 172 -349 178
rect -441 138 -412 172
rect -378 138 -349 172
rect -441 132 -349 138
rect -283 172 -191 178
rect -283 138 -254 172
rect -220 138 -191 172
rect -283 132 -191 138
rect -125 172 -33 178
rect -125 138 -96 172
rect -62 138 -33 172
rect -125 132 -33 138
rect 33 172 125 178
rect 33 138 62 172
rect 96 138 125 172
rect 33 132 125 138
rect 191 172 283 178
rect 191 138 220 172
rect 254 138 283 172
rect 191 132 283 138
rect 349 172 441 178
rect 349 138 378 172
rect 412 138 441 172
rect 349 132 441 138
rect 507 172 599 178
rect 507 138 536 172
rect 570 138 599 172
rect 507 132 599 138
rect 665 172 757 178
rect 665 138 694 172
rect 728 138 757 172
rect 665 132 757 138
rect 823 172 915 178
rect 823 138 852 172
rect 886 138 915 172
rect 823 132 915 138
rect 981 172 1073 178
rect 981 138 1010 172
rect 1044 138 1073 172
rect 981 132 1073 138
rect 1139 172 1231 178
rect 1139 138 1168 172
rect 1202 138 1231 172
rect 1139 132 1231 138
rect 1297 172 1389 178
rect 1297 138 1326 172
rect 1360 138 1389 172
rect 1297 132 1389 138
rect 1455 172 1547 178
rect 1455 138 1484 172
rect 1518 138 1547 172
rect 1455 132 1547 138
rect 1613 172 1705 178
rect 1613 138 1642 172
rect 1676 138 1705 172
rect 1613 132 1705 138
rect 1771 172 1863 178
rect 1771 138 1800 172
rect 1834 138 1863 172
rect 1771 132 1863 138
rect 1929 172 2021 178
rect 1929 138 1958 172
rect 1992 138 2021 172
rect 1929 132 2021 138
rect 2087 172 2179 178
rect 2087 138 2116 172
rect 2150 138 2179 172
rect 2087 132 2179 138
rect 2245 172 2337 178
rect 2245 138 2274 172
rect 2308 138 2337 172
rect 2245 132 2337 138
rect 2403 172 2495 178
rect 2403 138 2432 172
rect 2466 138 2495 172
rect 2403 132 2495 138
rect 2561 172 2653 178
rect 2561 138 2590 172
rect 2624 138 2653 172
rect 2561 132 2653 138
rect 2719 172 2811 178
rect 2719 138 2748 172
rect 2782 138 2811 172
rect 2719 132 2811 138
rect 2877 172 2969 178
rect 2877 138 2906 172
rect 2940 138 2969 172
rect 2877 132 2969 138
rect 3035 172 3127 178
rect 3035 138 3064 172
rect 3098 138 3127 172
rect 3035 132 3127 138
rect -3183 53 -3137 100
rect -3183 19 -3177 53
rect -3143 19 -3137 53
rect -3183 -19 -3137 19
rect -3183 -53 -3177 -19
rect -3143 -53 -3137 -19
rect -3183 -100 -3137 -53
rect -3025 53 -2979 100
rect -3025 19 -3019 53
rect -2985 19 -2979 53
rect -3025 -19 -2979 19
rect -3025 -53 -3019 -19
rect -2985 -53 -2979 -19
rect -3025 -100 -2979 -53
rect -2867 53 -2821 100
rect -2867 19 -2861 53
rect -2827 19 -2821 53
rect -2867 -19 -2821 19
rect -2867 -53 -2861 -19
rect -2827 -53 -2821 -19
rect -2867 -100 -2821 -53
rect -2709 53 -2663 100
rect -2709 19 -2703 53
rect -2669 19 -2663 53
rect -2709 -19 -2663 19
rect -2709 -53 -2703 -19
rect -2669 -53 -2663 -19
rect -2709 -100 -2663 -53
rect -2551 53 -2505 100
rect -2551 19 -2545 53
rect -2511 19 -2505 53
rect -2551 -19 -2505 19
rect -2551 -53 -2545 -19
rect -2511 -53 -2505 -19
rect -2551 -100 -2505 -53
rect -2393 53 -2347 100
rect -2393 19 -2387 53
rect -2353 19 -2347 53
rect -2393 -19 -2347 19
rect -2393 -53 -2387 -19
rect -2353 -53 -2347 -19
rect -2393 -100 -2347 -53
rect -2235 53 -2189 100
rect -2235 19 -2229 53
rect -2195 19 -2189 53
rect -2235 -19 -2189 19
rect -2235 -53 -2229 -19
rect -2195 -53 -2189 -19
rect -2235 -100 -2189 -53
rect -2077 53 -2031 100
rect -2077 19 -2071 53
rect -2037 19 -2031 53
rect -2077 -19 -2031 19
rect -2077 -53 -2071 -19
rect -2037 -53 -2031 -19
rect -2077 -100 -2031 -53
rect -1919 53 -1873 100
rect -1919 19 -1913 53
rect -1879 19 -1873 53
rect -1919 -19 -1873 19
rect -1919 -53 -1913 -19
rect -1879 -53 -1873 -19
rect -1919 -100 -1873 -53
rect -1761 53 -1715 100
rect -1761 19 -1755 53
rect -1721 19 -1715 53
rect -1761 -19 -1715 19
rect -1761 -53 -1755 -19
rect -1721 -53 -1715 -19
rect -1761 -100 -1715 -53
rect -1603 53 -1557 100
rect -1603 19 -1597 53
rect -1563 19 -1557 53
rect -1603 -19 -1557 19
rect -1603 -53 -1597 -19
rect -1563 -53 -1557 -19
rect -1603 -100 -1557 -53
rect -1445 53 -1399 100
rect -1445 19 -1439 53
rect -1405 19 -1399 53
rect -1445 -19 -1399 19
rect -1445 -53 -1439 -19
rect -1405 -53 -1399 -19
rect -1445 -100 -1399 -53
rect -1287 53 -1241 100
rect -1287 19 -1281 53
rect -1247 19 -1241 53
rect -1287 -19 -1241 19
rect -1287 -53 -1281 -19
rect -1247 -53 -1241 -19
rect -1287 -100 -1241 -53
rect -1129 53 -1083 100
rect -1129 19 -1123 53
rect -1089 19 -1083 53
rect -1129 -19 -1083 19
rect -1129 -53 -1123 -19
rect -1089 -53 -1083 -19
rect -1129 -100 -1083 -53
rect -971 53 -925 100
rect -971 19 -965 53
rect -931 19 -925 53
rect -971 -19 -925 19
rect -971 -53 -965 -19
rect -931 -53 -925 -19
rect -971 -100 -925 -53
rect -813 53 -767 100
rect -813 19 -807 53
rect -773 19 -767 53
rect -813 -19 -767 19
rect -813 -53 -807 -19
rect -773 -53 -767 -19
rect -813 -100 -767 -53
rect -655 53 -609 100
rect -655 19 -649 53
rect -615 19 -609 53
rect -655 -19 -609 19
rect -655 -53 -649 -19
rect -615 -53 -609 -19
rect -655 -100 -609 -53
rect -497 53 -451 100
rect -497 19 -491 53
rect -457 19 -451 53
rect -497 -19 -451 19
rect -497 -53 -491 -19
rect -457 -53 -451 -19
rect -497 -100 -451 -53
rect -339 53 -293 100
rect -339 19 -333 53
rect -299 19 -293 53
rect -339 -19 -293 19
rect -339 -53 -333 -19
rect -299 -53 -293 -19
rect -339 -100 -293 -53
rect -181 53 -135 100
rect -181 19 -175 53
rect -141 19 -135 53
rect -181 -19 -135 19
rect -181 -53 -175 -19
rect -141 -53 -135 -19
rect -181 -100 -135 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 135 53 181 100
rect 135 19 141 53
rect 175 19 181 53
rect 135 -19 181 19
rect 135 -53 141 -19
rect 175 -53 181 -19
rect 135 -100 181 -53
rect 293 53 339 100
rect 293 19 299 53
rect 333 19 339 53
rect 293 -19 339 19
rect 293 -53 299 -19
rect 333 -53 339 -19
rect 293 -100 339 -53
rect 451 53 497 100
rect 451 19 457 53
rect 491 19 497 53
rect 451 -19 497 19
rect 451 -53 457 -19
rect 491 -53 497 -19
rect 451 -100 497 -53
rect 609 53 655 100
rect 609 19 615 53
rect 649 19 655 53
rect 609 -19 655 19
rect 609 -53 615 -19
rect 649 -53 655 -19
rect 609 -100 655 -53
rect 767 53 813 100
rect 767 19 773 53
rect 807 19 813 53
rect 767 -19 813 19
rect 767 -53 773 -19
rect 807 -53 813 -19
rect 767 -100 813 -53
rect 925 53 971 100
rect 925 19 931 53
rect 965 19 971 53
rect 925 -19 971 19
rect 925 -53 931 -19
rect 965 -53 971 -19
rect 925 -100 971 -53
rect 1083 53 1129 100
rect 1083 19 1089 53
rect 1123 19 1129 53
rect 1083 -19 1129 19
rect 1083 -53 1089 -19
rect 1123 -53 1129 -19
rect 1083 -100 1129 -53
rect 1241 53 1287 100
rect 1241 19 1247 53
rect 1281 19 1287 53
rect 1241 -19 1287 19
rect 1241 -53 1247 -19
rect 1281 -53 1287 -19
rect 1241 -100 1287 -53
rect 1399 53 1445 100
rect 1399 19 1405 53
rect 1439 19 1445 53
rect 1399 -19 1445 19
rect 1399 -53 1405 -19
rect 1439 -53 1445 -19
rect 1399 -100 1445 -53
rect 1557 53 1603 100
rect 1557 19 1563 53
rect 1597 19 1603 53
rect 1557 -19 1603 19
rect 1557 -53 1563 -19
rect 1597 -53 1603 -19
rect 1557 -100 1603 -53
rect 1715 53 1761 100
rect 1715 19 1721 53
rect 1755 19 1761 53
rect 1715 -19 1761 19
rect 1715 -53 1721 -19
rect 1755 -53 1761 -19
rect 1715 -100 1761 -53
rect 1873 53 1919 100
rect 1873 19 1879 53
rect 1913 19 1919 53
rect 1873 -19 1919 19
rect 1873 -53 1879 -19
rect 1913 -53 1919 -19
rect 1873 -100 1919 -53
rect 2031 53 2077 100
rect 2031 19 2037 53
rect 2071 19 2077 53
rect 2031 -19 2077 19
rect 2031 -53 2037 -19
rect 2071 -53 2077 -19
rect 2031 -100 2077 -53
rect 2189 53 2235 100
rect 2189 19 2195 53
rect 2229 19 2235 53
rect 2189 -19 2235 19
rect 2189 -53 2195 -19
rect 2229 -53 2235 -19
rect 2189 -100 2235 -53
rect 2347 53 2393 100
rect 2347 19 2353 53
rect 2387 19 2393 53
rect 2347 -19 2393 19
rect 2347 -53 2353 -19
rect 2387 -53 2393 -19
rect 2347 -100 2393 -53
rect 2505 53 2551 100
rect 2505 19 2511 53
rect 2545 19 2551 53
rect 2505 -19 2551 19
rect 2505 -53 2511 -19
rect 2545 -53 2551 -19
rect 2505 -100 2551 -53
rect 2663 53 2709 100
rect 2663 19 2669 53
rect 2703 19 2709 53
rect 2663 -19 2709 19
rect 2663 -53 2669 -19
rect 2703 -53 2709 -19
rect 2663 -100 2709 -53
rect 2821 53 2867 100
rect 2821 19 2827 53
rect 2861 19 2867 53
rect 2821 -19 2867 19
rect 2821 -53 2827 -19
rect 2861 -53 2867 -19
rect 2821 -100 2867 -53
rect 2979 53 3025 100
rect 2979 19 2985 53
rect 3019 19 3025 53
rect 2979 -19 3025 19
rect 2979 -53 2985 -19
rect 3019 -53 3025 -19
rect 2979 -100 3025 -53
rect 3137 53 3183 100
rect 3137 19 3143 53
rect 3177 19 3183 53
rect 3137 -19 3183 19
rect 3137 -53 3143 -19
rect 3177 -53 3183 -19
rect 3137 -100 3183 -53
rect -3127 -138 -3035 -132
rect -3127 -172 -3098 -138
rect -3064 -172 -3035 -138
rect -3127 -178 -3035 -172
rect -2969 -138 -2877 -132
rect -2969 -172 -2940 -138
rect -2906 -172 -2877 -138
rect -2969 -178 -2877 -172
rect -2811 -138 -2719 -132
rect -2811 -172 -2782 -138
rect -2748 -172 -2719 -138
rect -2811 -178 -2719 -172
rect -2653 -138 -2561 -132
rect -2653 -172 -2624 -138
rect -2590 -172 -2561 -138
rect -2653 -178 -2561 -172
rect -2495 -138 -2403 -132
rect -2495 -172 -2466 -138
rect -2432 -172 -2403 -138
rect -2495 -178 -2403 -172
rect -2337 -138 -2245 -132
rect -2337 -172 -2308 -138
rect -2274 -172 -2245 -138
rect -2337 -178 -2245 -172
rect -2179 -138 -2087 -132
rect -2179 -172 -2150 -138
rect -2116 -172 -2087 -138
rect -2179 -178 -2087 -172
rect -2021 -138 -1929 -132
rect -2021 -172 -1992 -138
rect -1958 -172 -1929 -138
rect -2021 -178 -1929 -172
rect -1863 -138 -1771 -132
rect -1863 -172 -1834 -138
rect -1800 -172 -1771 -138
rect -1863 -178 -1771 -172
rect -1705 -138 -1613 -132
rect -1705 -172 -1676 -138
rect -1642 -172 -1613 -138
rect -1705 -178 -1613 -172
rect -1547 -138 -1455 -132
rect -1547 -172 -1518 -138
rect -1484 -172 -1455 -138
rect -1547 -178 -1455 -172
rect -1389 -138 -1297 -132
rect -1389 -172 -1360 -138
rect -1326 -172 -1297 -138
rect -1389 -178 -1297 -172
rect -1231 -138 -1139 -132
rect -1231 -172 -1202 -138
rect -1168 -172 -1139 -138
rect -1231 -178 -1139 -172
rect -1073 -138 -981 -132
rect -1073 -172 -1044 -138
rect -1010 -172 -981 -138
rect -1073 -178 -981 -172
rect -915 -138 -823 -132
rect -915 -172 -886 -138
rect -852 -172 -823 -138
rect -915 -178 -823 -172
rect -757 -138 -665 -132
rect -757 -172 -728 -138
rect -694 -172 -665 -138
rect -757 -178 -665 -172
rect -599 -138 -507 -132
rect -599 -172 -570 -138
rect -536 -172 -507 -138
rect -599 -178 -507 -172
rect -441 -138 -349 -132
rect -441 -172 -412 -138
rect -378 -172 -349 -138
rect -441 -178 -349 -172
rect -283 -138 -191 -132
rect -283 -172 -254 -138
rect -220 -172 -191 -138
rect -283 -178 -191 -172
rect -125 -138 -33 -132
rect -125 -172 -96 -138
rect -62 -172 -33 -138
rect -125 -178 -33 -172
rect 33 -138 125 -132
rect 33 -172 62 -138
rect 96 -172 125 -138
rect 33 -178 125 -172
rect 191 -138 283 -132
rect 191 -172 220 -138
rect 254 -172 283 -138
rect 191 -178 283 -172
rect 349 -138 441 -132
rect 349 -172 378 -138
rect 412 -172 441 -138
rect 349 -178 441 -172
rect 507 -138 599 -132
rect 507 -172 536 -138
rect 570 -172 599 -138
rect 507 -178 599 -172
rect 665 -138 757 -132
rect 665 -172 694 -138
rect 728 -172 757 -138
rect 665 -178 757 -172
rect 823 -138 915 -132
rect 823 -172 852 -138
rect 886 -172 915 -138
rect 823 -178 915 -172
rect 981 -138 1073 -132
rect 981 -172 1010 -138
rect 1044 -172 1073 -138
rect 981 -178 1073 -172
rect 1139 -138 1231 -132
rect 1139 -172 1168 -138
rect 1202 -172 1231 -138
rect 1139 -178 1231 -172
rect 1297 -138 1389 -132
rect 1297 -172 1326 -138
rect 1360 -172 1389 -138
rect 1297 -178 1389 -172
rect 1455 -138 1547 -132
rect 1455 -172 1484 -138
rect 1518 -172 1547 -138
rect 1455 -178 1547 -172
rect 1613 -138 1705 -132
rect 1613 -172 1642 -138
rect 1676 -172 1705 -138
rect 1613 -178 1705 -172
rect 1771 -138 1863 -132
rect 1771 -172 1800 -138
rect 1834 -172 1863 -138
rect 1771 -178 1863 -172
rect 1929 -138 2021 -132
rect 1929 -172 1958 -138
rect 1992 -172 2021 -138
rect 1929 -178 2021 -172
rect 2087 -138 2179 -132
rect 2087 -172 2116 -138
rect 2150 -172 2179 -138
rect 2087 -178 2179 -172
rect 2245 -138 2337 -132
rect 2245 -172 2274 -138
rect 2308 -172 2337 -138
rect 2245 -178 2337 -172
rect 2403 -138 2495 -132
rect 2403 -172 2432 -138
rect 2466 -172 2495 -138
rect 2403 -178 2495 -172
rect 2561 -138 2653 -132
rect 2561 -172 2590 -138
rect 2624 -172 2653 -138
rect 2561 -178 2653 -172
rect 2719 -138 2811 -132
rect 2719 -172 2748 -138
rect 2782 -172 2811 -138
rect 2719 -178 2811 -172
rect 2877 -138 2969 -132
rect 2877 -172 2906 -138
rect 2940 -172 2969 -138
rect 2877 -178 2969 -172
rect 3035 -138 3127 -132
rect 3035 -172 3064 -138
rect 3098 -172 3127 -138
rect 3035 -178 3127 -172
rect -3127 -246 -3035 -240
rect -3127 -280 -3098 -246
rect -3064 -280 -3035 -246
rect -3127 -286 -3035 -280
rect -2969 -246 -2877 -240
rect -2969 -280 -2940 -246
rect -2906 -280 -2877 -246
rect -2969 -286 -2877 -280
rect -2811 -246 -2719 -240
rect -2811 -280 -2782 -246
rect -2748 -280 -2719 -246
rect -2811 -286 -2719 -280
rect -2653 -246 -2561 -240
rect -2653 -280 -2624 -246
rect -2590 -280 -2561 -246
rect -2653 -286 -2561 -280
rect -2495 -246 -2403 -240
rect -2495 -280 -2466 -246
rect -2432 -280 -2403 -246
rect -2495 -286 -2403 -280
rect -2337 -246 -2245 -240
rect -2337 -280 -2308 -246
rect -2274 -280 -2245 -246
rect -2337 -286 -2245 -280
rect -2179 -246 -2087 -240
rect -2179 -280 -2150 -246
rect -2116 -280 -2087 -246
rect -2179 -286 -2087 -280
rect -2021 -246 -1929 -240
rect -2021 -280 -1992 -246
rect -1958 -280 -1929 -246
rect -2021 -286 -1929 -280
rect -1863 -246 -1771 -240
rect -1863 -280 -1834 -246
rect -1800 -280 -1771 -246
rect -1863 -286 -1771 -280
rect -1705 -246 -1613 -240
rect -1705 -280 -1676 -246
rect -1642 -280 -1613 -246
rect -1705 -286 -1613 -280
rect -1547 -246 -1455 -240
rect -1547 -280 -1518 -246
rect -1484 -280 -1455 -246
rect -1547 -286 -1455 -280
rect -1389 -246 -1297 -240
rect -1389 -280 -1360 -246
rect -1326 -280 -1297 -246
rect -1389 -286 -1297 -280
rect -1231 -246 -1139 -240
rect -1231 -280 -1202 -246
rect -1168 -280 -1139 -246
rect -1231 -286 -1139 -280
rect -1073 -246 -981 -240
rect -1073 -280 -1044 -246
rect -1010 -280 -981 -246
rect -1073 -286 -981 -280
rect -915 -246 -823 -240
rect -915 -280 -886 -246
rect -852 -280 -823 -246
rect -915 -286 -823 -280
rect -757 -246 -665 -240
rect -757 -280 -728 -246
rect -694 -280 -665 -246
rect -757 -286 -665 -280
rect -599 -246 -507 -240
rect -599 -280 -570 -246
rect -536 -280 -507 -246
rect -599 -286 -507 -280
rect -441 -246 -349 -240
rect -441 -280 -412 -246
rect -378 -280 -349 -246
rect -441 -286 -349 -280
rect -283 -246 -191 -240
rect -283 -280 -254 -246
rect -220 -280 -191 -246
rect -283 -286 -191 -280
rect -125 -246 -33 -240
rect -125 -280 -96 -246
rect -62 -280 -33 -246
rect -125 -286 -33 -280
rect 33 -246 125 -240
rect 33 -280 62 -246
rect 96 -280 125 -246
rect 33 -286 125 -280
rect 191 -246 283 -240
rect 191 -280 220 -246
rect 254 -280 283 -246
rect 191 -286 283 -280
rect 349 -246 441 -240
rect 349 -280 378 -246
rect 412 -280 441 -246
rect 349 -286 441 -280
rect 507 -246 599 -240
rect 507 -280 536 -246
rect 570 -280 599 -246
rect 507 -286 599 -280
rect 665 -246 757 -240
rect 665 -280 694 -246
rect 728 -280 757 -246
rect 665 -286 757 -280
rect 823 -246 915 -240
rect 823 -280 852 -246
rect 886 -280 915 -246
rect 823 -286 915 -280
rect 981 -246 1073 -240
rect 981 -280 1010 -246
rect 1044 -280 1073 -246
rect 981 -286 1073 -280
rect 1139 -246 1231 -240
rect 1139 -280 1168 -246
rect 1202 -280 1231 -246
rect 1139 -286 1231 -280
rect 1297 -246 1389 -240
rect 1297 -280 1326 -246
rect 1360 -280 1389 -246
rect 1297 -286 1389 -280
rect 1455 -246 1547 -240
rect 1455 -280 1484 -246
rect 1518 -280 1547 -246
rect 1455 -286 1547 -280
rect 1613 -246 1705 -240
rect 1613 -280 1642 -246
rect 1676 -280 1705 -246
rect 1613 -286 1705 -280
rect 1771 -246 1863 -240
rect 1771 -280 1800 -246
rect 1834 -280 1863 -246
rect 1771 -286 1863 -280
rect 1929 -246 2021 -240
rect 1929 -280 1958 -246
rect 1992 -280 2021 -246
rect 1929 -286 2021 -280
rect 2087 -246 2179 -240
rect 2087 -280 2116 -246
rect 2150 -280 2179 -246
rect 2087 -286 2179 -280
rect 2245 -246 2337 -240
rect 2245 -280 2274 -246
rect 2308 -280 2337 -246
rect 2245 -286 2337 -280
rect 2403 -246 2495 -240
rect 2403 -280 2432 -246
rect 2466 -280 2495 -246
rect 2403 -286 2495 -280
rect 2561 -246 2653 -240
rect 2561 -280 2590 -246
rect 2624 -280 2653 -246
rect 2561 -286 2653 -280
rect 2719 -246 2811 -240
rect 2719 -280 2748 -246
rect 2782 -280 2811 -246
rect 2719 -286 2811 -280
rect 2877 -246 2969 -240
rect 2877 -280 2906 -246
rect 2940 -280 2969 -246
rect 2877 -286 2969 -280
rect 3035 -246 3127 -240
rect 3035 -280 3064 -246
rect 3098 -280 3127 -246
rect 3035 -286 3127 -280
rect -3183 -365 -3137 -318
rect -3183 -399 -3177 -365
rect -3143 -399 -3137 -365
rect -3183 -437 -3137 -399
rect -3183 -471 -3177 -437
rect -3143 -471 -3137 -437
rect -3183 -518 -3137 -471
rect -3025 -365 -2979 -318
rect -3025 -399 -3019 -365
rect -2985 -399 -2979 -365
rect -3025 -437 -2979 -399
rect -3025 -471 -3019 -437
rect -2985 -471 -2979 -437
rect -3025 -518 -2979 -471
rect -2867 -365 -2821 -318
rect -2867 -399 -2861 -365
rect -2827 -399 -2821 -365
rect -2867 -437 -2821 -399
rect -2867 -471 -2861 -437
rect -2827 -471 -2821 -437
rect -2867 -518 -2821 -471
rect -2709 -365 -2663 -318
rect -2709 -399 -2703 -365
rect -2669 -399 -2663 -365
rect -2709 -437 -2663 -399
rect -2709 -471 -2703 -437
rect -2669 -471 -2663 -437
rect -2709 -518 -2663 -471
rect -2551 -365 -2505 -318
rect -2551 -399 -2545 -365
rect -2511 -399 -2505 -365
rect -2551 -437 -2505 -399
rect -2551 -471 -2545 -437
rect -2511 -471 -2505 -437
rect -2551 -518 -2505 -471
rect -2393 -365 -2347 -318
rect -2393 -399 -2387 -365
rect -2353 -399 -2347 -365
rect -2393 -437 -2347 -399
rect -2393 -471 -2387 -437
rect -2353 -471 -2347 -437
rect -2393 -518 -2347 -471
rect -2235 -365 -2189 -318
rect -2235 -399 -2229 -365
rect -2195 -399 -2189 -365
rect -2235 -437 -2189 -399
rect -2235 -471 -2229 -437
rect -2195 -471 -2189 -437
rect -2235 -518 -2189 -471
rect -2077 -365 -2031 -318
rect -2077 -399 -2071 -365
rect -2037 -399 -2031 -365
rect -2077 -437 -2031 -399
rect -2077 -471 -2071 -437
rect -2037 -471 -2031 -437
rect -2077 -518 -2031 -471
rect -1919 -365 -1873 -318
rect -1919 -399 -1913 -365
rect -1879 -399 -1873 -365
rect -1919 -437 -1873 -399
rect -1919 -471 -1913 -437
rect -1879 -471 -1873 -437
rect -1919 -518 -1873 -471
rect -1761 -365 -1715 -318
rect -1761 -399 -1755 -365
rect -1721 -399 -1715 -365
rect -1761 -437 -1715 -399
rect -1761 -471 -1755 -437
rect -1721 -471 -1715 -437
rect -1761 -518 -1715 -471
rect -1603 -365 -1557 -318
rect -1603 -399 -1597 -365
rect -1563 -399 -1557 -365
rect -1603 -437 -1557 -399
rect -1603 -471 -1597 -437
rect -1563 -471 -1557 -437
rect -1603 -518 -1557 -471
rect -1445 -365 -1399 -318
rect -1445 -399 -1439 -365
rect -1405 -399 -1399 -365
rect -1445 -437 -1399 -399
rect -1445 -471 -1439 -437
rect -1405 -471 -1399 -437
rect -1445 -518 -1399 -471
rect -1287 -365 -1241 -318
rect -1287 -399 -1281 -365
rect -1247 -399 -1241 -365
rect -1287 -437 -1241 -399
rect -1287 -471 -1281 -437
rect -1247 -471 -1241 -437
rect -1287 -518 -1241 -471
rect -1129 -365 -1083 -318
rect -1129 -399 -1123 -365
rect -1089 -399 -1083 -365
rect -1129 -437 -1083 -399
rect -1129 -471 -1123 -437
rect -1089 -471 -1083 -437
rect -1129 -518 -1083 -471
rect -971 -365 -925 -318
rect -971 -399 -965 -365
rect -931 -399 -925 -365
rect -971 -437 -925 -399
rect -971 -471 -965 -437
rect -931 -471 -925 -437
rect -971 -518 -925 -471
rect -813 -365 -767 -318
rect -813 -399 -807 -365
rect -773 -399 -767 -365
rect -813 -437 -767 -399
rect -813 -471 -807 -437
rect -773 -471 -767 -437
rect -813 -518 -767 -471
rect -655 -365 -609 -318
rect -655 -399 -649 -365
rect -615 -399 -609 -365
rect -655 -437 -609 -399
rect -655 -471 -649 -437
rect -615 -471 -609 -437
rect -655 -518 -609 -471
rect -497 -365 -451 -318
rect -497 -399 -491 -365
rect -457 -399 -451 -365
rect -497 -437 -451 -399
rect -497 -471 -491 -437
rect -457 -471 -451 -437
rect -497 -518 -451 -471
rect -339 -365 -293 -318
rect -339 -399 -333 -365
rect -299 -399 -293 -365
rect -339 -437 -293 -399
rect -339 -471 -333 -437
rect -299 -471 -293 -437
rect -339 -518 -293 -471
rect -181 -365 -135 -318
rect -181 -399 -175 -365
rect -141 -399 -135 -365
rect -181 -437 -135 -399
rect -181 -471 -175 -437
rect -141 -471 -135 -437
rect -181 -518 -135 -471
rect -23 -365 23 -318
rect -23 -399 -17 -365
rect 17 -399 23 -365
rect -23 -437 23 -399
rect -23 -471 -17 -437
rect 17 -471 23 -437
rect -23 -518 23 -471
rect 135 -365 181 -318
rect 135 -399 141 -365
rect 175 -399 181 -365
rect 135 -437 181 -399
rect 135 -471 141 -437
rect 175 -471 181 -437
rect 135 -518 181 -471
rect 293 -365 339 -318
rect 293 -399 299 -365
rect 333 -399 339 -365
rect 293 -437 339 -399
rect 293 -471 299 -437
rect 333 -471 339 -437
rect 293 -518 339 -471
rect 451 -365 497 -318
rect 451 -399 457 -365
rect 491 -399 497 -365
rect 451 -437 497 -399
rect 451 -471 457 -437
rect 491 -471 497 -437
rect 451 -518 497 -471
rect 609 -365 655 -318
rect 609 -399 615 -365
rect 649 -399 655 -365
rect 609 -437 655 -399
rect 609 -471 615 -437
rect 649 -471 655 -437
rect 609 -518 655 -471
rect 767 -365 813 -318
rect 767 -399 773 -365
rect 807 -399 813 -365
rect 767 -437 813 -399
rect 767 -471 773 -437
rect 807 -471 813 -437
rect 767 -518 813 -471
rect 925 -365 971 -318
rect 925 -399 931 -365
rect 965 -399 971 -365
rect 925 -437 971 -399
rect 925 -471 931 -437
rect 965 -471 971 -437
rect 925 -518 971 -471
rect 1083 -365 1129 -318
rect 1083 -399 1089 -365
rect 1123 -399 1129 -365
rect 1083 -437 1129 -399
rect 1083 -471 1089 -437
rect 1123 -471 1129 -437
rect 1083 -518 1129 -471
rect 1241 -365 1287 -318
rect 1241 -399 1247 -365
rect 1281 -399 1287 -365
rect 1241 -437 1287 -399
rect 1241 -471 1247 -437
rect 1281 -471 1287 -437
rect 1241 -518 1287 -471
rect 1399 -365 1445 -318
rect 1399 -399 1405 -365
rect 1439 -399 1445 -365
rect 1399 -437 1445 -399
rect 1399 -471 1405 -437
rect 1439 -471 1445 -437
rect 1399 -518 1445 -471
rect 1557 -365 1603 -318
rect 1557 -399 1563 -365
rect 1597 -399 1603 -365
rect 1557 -437 1603 -399
rect 1557 -471 1563 -437
rect 1597 -471 1603 -437
rect 1557 -518 1603 -471
rect 1715 -365 1761 -318
rect 1715 -399 1721 -365
rect 1755 -399 1761 -365
rect 1715 -437 1761 -399
rect 1715 -471 1721 -437
rect 1755 -471 1761 -437
rect 1715 -518 1761 -471
rect 1873 -365 1919 -318
rect 1873 -399 1879 -365
rect 1913 -399 1919 -365
rect 1873 -437 1919 -399
rect 1873 -471 1879 -437
rect 1913 -471 1919 -437
rect 1873 -518 1919 -471
rect 2031 -365 2077 -318
rect 2031 -399 2037 -365
rect 2071 -399 2077 -365
rect 2031 -437 2077 -399
rect 2031 -471 2037 -437
rect 2071 -471 2077 -437
rect 2031 -518 2077 -471
rect 2189 -365 2235 -318
rect 2189 -399 2195 -365
rect 2229 -399 2235 -365
rect 2189 -437 2235 -399
rect 2189 -471 2195 -437
rect 2229 -471 2235 -437
rect 2189 -518 2235 -471
rect 2347 -365 2393 -318
rect 2347 -399 2353 -365
rect 2387 -399 2393 -365
rect 2347 -437 2393 -399
rect 2347 -471 2353 -437
rect 2387 -471 2393 -437
rect 2347 -518 2393 -471
rect 2505 -365 2551 -318
rect 2505 -399 2511 -365
rect 2545 -399 2551 -365
rect 2505 -437 2551 -399
rect 2505 -471 2511 -437
rect 2545 -471 2551 -437
rect 2505 -518 2551 -471
rect 2663 -365 2709 -318
rect 2663 -399 2669 -365
rect 2703 -399 2709 -365
rect 2663 -437 2709 -399
rect 2663 -471 2669 -437
rect 2703 -471 2709 -437
rect 2663 -518 2709 -471
rect 2821 -365 2867 -318
rect 2821 -399 2827 -365
rect 2861 -399 2867 -365
rect 2821 -437 2867 -399
rect 2821 -471 2827 -437
rect 2861 -471 2867 -437
rect 2821 -518 2867 -471
rect 2979 -365 3025 -318
rect 2979 -399 2985 -365
rect 3019 -399 3025 -365
rect 2979 -437 3025 -399
rect 2979 -471 2985 -437
rect 3019 -471 3025 -437
rect 2979 -518 3025 -471
rect 3137 -365 3183 -318
rect 3137 -399 3143 -365
rect 3177 -399 3183 -365
rect 3137 -437 3183 -399
rect 3137 -471 3143 -437
rect 3177 -471 3183 -437
rect 3137 -518 3183 -471
rect -3127 -556 -3035 -550
rect -3127 -590 -3098 -556
rect -3064 -590 -3035 -556
rect -3127 -596 -3035 -590
rect -2969 -556 -2877 -550
rect -2969 -590 -2940 -556
rect -2906 -590 -2877 -556
rect -2969 -596 -2877 -590
rect -2811 -556 -2719 -550
rect -2811 -590 -2782 -556
rect -2748 -590 -2719 -556
rect -2811 -596 -2719 -590
rect -2653 -556 -2561 -550
rect -2653 -590 -2624 -556
rect -2590 -590 -2561 -556
rect -2653 -596 -2561 -590
rect -2495 -556 -2403 -550
rect -2495 -590 -2466 -556
rect -2432 -590 -2403 -556
rect -2495 -596 -2403 -590
rect -2337 -556 -2245 -550
rect -2337 -590 -2308 -556
rect -2274 -590 -2245 -556
rect -2337 -596 -2245 -590
rect -2179 -556 -2087 -550
rect -2179 -590 -2150 -556
rect -2116 -590 -2087 -556
rect -2179 -596 -2087 -590
rect -2021 -556 -1929 -550
rect -2021 -590 -1992 -556
rect -1958 -590 -1929 -556
rect -2021 -596 -1929 -590
rect -1863 -556 -1771 -550
rect -1863 -590 -1834 -556
rect -1800 -590 -1771 -556
rect -1863 -596 -1771 -590
rect -1705 -556 -1613 -550
rect -1705 -590 -1676 -556
rect -1642 -590 -1613 -556
rect -1705 -596 -1613 -590
rect -1547 -556 -1455 -550
rect -1547 -590 -1518 -556
rect -1484 -590 -1455 -556
rect -1547 -596 -1455 -590
rect -1389 -556 -1297 -550
rect -1389 -590 -1360 -556
rect -1326 -590 -1297 -556
rect -1389 -596 -1297 -590
rect -1231 -556 -1139 -550
rect -1231 -590 -1202 -556
rect -1168 -590 -1139 -556
rect -1231 -596 -1139 -590
rect -1073 -556 -981 -550
rect -1073 -590 -1044 -556
rect -1010 -590 -981 -556
rect -1073 -596 -981 -590
rect -915 -556 -823 -550
rect -915 -590 -886 -556
rect -852 -590 -823 -556
rect -915 -596 -823 -590
rect -757 -556 -665 -550
rect -757 -590 -728 -556
rect -694 -590 -665 -556
rect -757 -596 -665 -590
rect -599 -556 -507 -550
rect -599 -590 -570 -556
rect -536 -590 -507 -556
rect -599 -596 -507 -590
rect -441 -556 -349 -550
rect -441 -590 -412 -556
rect -378 -590 -349 -556
rect -441 -596 -349 -590
rect -283 -556 -191 -550
rect -283 -590 -254 -556
rect -220 -590 -191 -556
rect -283 -596 -191 -590
rect -125 -556 -33 -550
rect -125 -590 -96 -556
rect -62 -590 -33 -556
rect -125 -596 -33 -590
rect 33 -556 125 -550
rect 33 -590 62 -556
rect 96 -590 125 -556
rect 33 -596 125 -590
rect 191 -556 283 -550
rect 191 -590 220 -556
rect 254 -590 283 -556
rect 191 -596 283 -590
rect 349 -556 441 -550
rect 349 -590 378 -556
rect 412 -590 441 -556
rect 349 -596 441 -590
rect 507 -556 599 -550
rect 507 -590 536 -556
rect 570 -590 599 -556
rect 507 -596 599 -590
rect 665 -556 757 -550
rect 665 -590 694 -556
rect 728 -590 757 -556
rect 665 -596 757 -590
rect 823 -556 915 -550
rect 823 -590 852 -556
rect 886 -590 915 -556
rect 823 -596 915 -590
rect 981 -556 1073 -550
rect 981 -590 1010 -556
rect 1044 -590 1073 -556
rect 981 -596 1073 -590
rect 1139 -556 1231 -550
rect 1139 -590 1168 -556
rect 1202 -590 1231 -556
rect 1139 -596 1231 -590
rect 1297 -556 1389 -550
rect 1297 -590 1326 -556
rect 1360 -590 1389 -556
rect 1297 -596 1389 -590
rect 1455 -556 1547 -550
rect 1455 -590 1484 -556
rect 1518 -590 1547 -556
rect 1455 -596 1547 -590
rect 1613 -556 1705 -550
rect 1613 -590 1642 -556
rect 1676 -590 1705 -556
rect 1613 -596 1705 -590
rect 1771 -556 1863 -550
rect 1771 -590 1800 -556
rect 1834 -590 1863 -556
rect 1771 -596 1863 -590
rect 1929 -556 2021 -550
rect 1929 -590 1958 -556
rect 1992 -590 2021 -556
rect 1929 -596 2021 -590
rect 2087 -556 2179 -550
rect 2087 -590 2116 -556
rect 2150 -590 2179 -556
rect 2087 -596 2179 -590
rect 2245 -556 2337 -550
rect 2245 -590 2274 -556
rect 2308 -590 2337 -556
rect 2245 -596 2337 -590
rect 2403 -556 2495 -550
rect 2403 -590 2432 -556
rect 2466 -590 2495 -556
rect 2403 -596 2495 -590
rect 2561 -556 2653 -550
rect 2561 -590 2590 -556
rect 2624 -590 2653 -556
rect 2561 -596 2653 -590
rect 2719 -556 2811 -550
rect 2719 -590 2748 -556
rect 2782 -590 2811 -556
rect 2719 -596 2811 -590
rect 2877 -556 2969 -550
rect 2877 -590 2906 -556
rect 2940 -590 2969 -556
rect 2877 -596 2969 -590
rect 3035 -556 3127 -550
rect 3035 -590 3064 -556
rect 3098 -590 3127 -556
rect 3035 -596 3127 -590
<< properties >>
string FIXED_BBOX -3294 -711 3294 711
<< end >>
