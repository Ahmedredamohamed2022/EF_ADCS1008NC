magic
tech sky130A
magscale 1 2
timestamp 1693827120
<< pwell >>
rect -505 -348 505 348
<< mvnmos >>
rect -287 -100 -187 100
rect -129 -100 -29 100
rect 29 -100 129 100
rect 187 -100 287 100
<< mvndiff >>
rect -345 85 -287 100
rect -345 51 -333 85
rect -299 51 -287 85
rect -345 17 -287 51
rect -345 -17 -333 17
rect -299 -17 -287 17
rect -345 -51 -287 -17
rect -345 -85 -333 -51
rect -299 -85 -287 -51
rect -345 -100 -287 -85
rect -187 85 -129 100
rect -187 51 -175 85
rect -141 51 -129 85
rect -187 17 -129 51
rect -187 -17 -175 17
rect -141 -17 -129 17
rect -187 -51 -129 -17
rect -187 -85 -175 -51
rect -141 -85 -129 -51
rect -187 -100 -129 -85
rect -29 85 29 100
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -100 29 -85
rect 129 85 187 100
rect 129 51 141 85
rect 175 51 187 85
rect 129 17 187 51
rect 129 -17 141 17
rect 175 -17 187 17
rect 129 -51 187 -17
rect 129 -85 141 -51
rect 175 -85 187 -51
rect 129 -100 187 -85
rect 287 85 345 100
rect 287 51 299 85
rect 333 51 345 85
rect 287 17 345 51
rect 287 -17 299 17
rect 333 -17 345 17
rect 287 -51 345 -17
rect 287 -85 299 -51
rect 333 -85 345 -51
rect 287 -100 345 -85
<< mvndiffc >>
rect -333 51 -299 85
rect -333 -17 -299 17
rect -333 -85 -299 -51
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect 299 51 333 85
rect 299 -17 333 17
rect 299 -85 333 -51
<< mvpsubdiff >>
rect -479 310 479 322
rect -479 276 -357 310
rect -323 276 -289 310
rect -255 276 -221 310
rect -187 276 -153 310
rect -119 276 -85 310
rect -51 276 -17 310
rect 17 276 51 310
rect 85 276 119 310
rect 153 276 187 310
rect 221 276 255 310
rect 289 276 323 310
rect 357 276 479 310
rect -479 264 479 276
rect -479 187 -421 264
rect -479 153 -467 187
rect -433 153 -421 187
rect -479 119 -421 153
rect -479 85 -467 119
rect -433 85 -421 119
rect 421 187 479 264
rect 421 153 433 187
rect 467 153 479 187
rect 421 119 479 153
rect -479 51 -421 85
rect -479 17 -467 51
rect -433 17 -421 51
rect -479 -17 -421 17
rect -479 -51 -467 -17
rect -433 -51 -421 -17
rect -479 -85 -421 -51
rect -479 -119 -467 -85
rect -433 -119 -421 -85
rect 421 85 433 119
rect 467 85 479 119
rect 421 51 479 85
rect 421 17 433 51
rect 467 17 479 51
rect 421 -17 479 17
rect 421 -51 433 -17
rect 467 -51 479 -17
rect 421 -85 479 -51
rect -479 -153 -421 -119
rect -479 -187 -467 -153
rect -433 -187 -421 -153
rect -479 -264 -421 -187
rect 421 -119 433 -85
rect 467 -119 479 -85
rect 421 -153 479 -119
rect 421 -187 433 -153
rect 467 -187 479 -153
rect 421 -264 479 -187
rect -479 -276 479 -264
rect -479 -310 -357 -276
rect -323 -310 -289 -276
rect -255 -310 -221 -276
rect -187 -310 -153 -276
rect -119 -310 -85 -276
rect -51 -310 -17 -276
rect 17 -310 51 -276
rect 85 -310 119 -276
rect 153 -310 187 -276
rect 221 -310 255 -276
rect 289 -310 323 -276
rect 357 -310 479 -276
rect -479 -322 479 -310
<< mvpsubdiffcont >>
rect -357 276 -323 310
rect -289 276 -255 310
rect -221 276 -187 310
rect -153 276 -119 310
rect -85 276 -51 310
rect -17 276 17 310
rect 51 276 85 310
rect 119 276 153 310
rect 187 276 221 310
rect 255 276 289 310
rect 323 276 357 310
rect -467 153 -433 187
rect -467 85 -433 119
rect 433 153 467 187
rect -467 17 -433 51
rect -467 -51 -433 -17
rect -467 -119 -433 -85
rect 433 85 467 119
rect 433 17 467 51
rect 433 -51 467 -17
rect -467 -187 -433 -153
rect 433 -119 467 -85
rect 433 -187 467 -153
rect -357 -310 -323 -276
rect -289 -310 -255 -276
rect -221 -310 -187 -276
rect -153 -310 -119 -276
rect -85 -310 -51 -276
rect -17 -310 17 -276
rect 51 -310 85 -276
rect 119 -310 153 -276
rect 187 -310 221 -276
rect 255 -310 289 -276
rect 323 -310 357 -276
<< poly >>
rect -287 172 -187 188
rect -287 138 -254 172
rect -220 138 -187 172
rect -287 100 -187 138
rect -129 172 -29 188
rect -129 138 -96 172
rect -62 138 -29 172
rect -129 100 -29 138
rect 29 172 129 188
rect 29 138 62 172
rect 96 138 129 172
rect 29 100 129 138
rect 187 172 287 188
rect 187 138 220 172
rect 254 138 287 172
rect 187 100 287 138
rect -287 -138 -187 -100
rect -287 -172 -254 -138
rect -220 -172 -187 -138
rect -287 -188 -187 -172
rect -129 -138 -29 -100
rect -129 -172 -96 -138
rect -62 -172 -29 -138
rect -129 -188 -29 -172
rect 29 -138 129 -100
rect 29 -172 62 -138
rect 96 -172 129 -138
rect 29 -188 129 -172
rect 187 -138 287 -100
rect 187 -172 220 -138
rect 254 -172 287 -138
rect 187 -188 287 -172
<< polycont >>
rect -254 138 -220 172
rect -96 138 -62 172
rect 62 138 96 172
rect 220 138 254 172
rect -254 -172 -220 -138
rect -96 -172 -62 -138
rect 62 -172 96 -138
rect 220 -172 254 -138
<< locali >>
rect -467 276 -357 310
rect -323 276 -289 310
rect -255 276 -221 310
rect -187 276 -153 310
rect -119 276 -85 310
rect -51 276 -17 310
rect 17 276 51 310
rect 85 276 119 310
rect 153 276 187 310
rect 221 276 255 310
rect 289 276 323 310
rect 357 276 467 310
rect -467 187 -433 276
rect 433 187 467 276
rect -467 119 -433 153
rect -287 138 -254 172
rect -220 138 -187 172
rect -129 138 -96 172
rect -62 138 -29 172
rect 29 138 62 172
rect 96 138 129 172
rect 187 138 220 172
rect 254 138 287 172
rect 433 119 467 153
rect -467 51 -433 85
rect -467 -17 -433 17
rect -467 -85 -433 -51
rect -333 85 -299 104
rect -333 17 -299 19
rect -333 -19 -299 -17
rect -333 -104 -299 -85
rect -175 85 -141 104
rect -175 17 -141 19
rect -175 -19 -141 -17
rect -175 -104 -141 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 141 85 175 104
rect 141 17 175 19
rect 141 -19 175 -17
rect 141 -104 175 -85
rect 299 85 333 104
rect 299 17 333 19
rect 299 -19 333 -17
rect 299 -104 333 -85
rect 433 51 467 85
rect 433 -17 467 17
rect 433 -85 467 -51
rect -467 -153 -433 -119
rect -287 -172 -254 -138
rect -220 -172 -187 -138
rect -129 -172 -96 -138
rect -62 -172 -29 -138
rect 29 -172 62 -138
rect 96 -172 129 -138
rect 187 -172 220 -138
rect 254 -172 287 -138
rect 433 -153 467 -119
rect -467 -276 -433 -187
rect 433 -276 467 -187
rect -467 -310 -357 -276
rect -323 -310 -289 -276
rect -255 -310 -221 -276
rect -187 -310 -153 -276
rect -119 -310 -85 -276
rect -51 -310 -17 -276
rect 17 -310 51 -276
rect 85 -310 119 -276
rect 153 -310 187 -276
rect 221 -310 255 -276
rect 289 -310 323 -276
rect 357 -310 467 -276
<< viali >>
rect -254 138 -220 172
rect -96 138 -62 172
rect 62 138 96 172
rect 220 138 254 172
rect -333 51 -299 53
rect -333 19 -299 51
rect -333 -51 -299 -19
rect -333 -53 -299 -51
rect -175 51 -141 53
rect -175 19 -141 51
rect -175 -51 -141 -19
rect -175 -53 -141 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 141 51 175 53
rect 141 19 175 51
rect 141 -51 175 -19
rect 141 -53 175 -51
rect 299 51 333 53
rect 299 19 333 51
rect 299 -51 333 -19
rect 299 -53 333 -51
rect -254 -172 -220 -138
rect -96 -172 -62 -138
rect 62 -172 96 -138
rect 220 -172 254 -138
<< metal1 >>
rect -283 172 -191 178
rect -283 138 -254 172
rect -220 138 -191 172
rect -283 132 -191 138
rect -125 172 -33 178
rect -125 138 -96 172
rect -62 138 -33 172
rect -125 132 -33 138
rect 33 172 125 178
rect 33 138 62 172
rect 96 138 125 172
rect 33 132 125 138
rect 191 172 283 178
rect 191 138 220 172
rect 254 138 283 172
rect 191 132 283 138
rect -339 53 -293 100
rect -339 19 -333 53
rect -299 19 -293 53
rect -339 -19 -293 19
rect -339 -53 -333 -19
rect -299 -53 -293 -19
rect -339 -100 -293 -53
rect -181 53 -135 100
rect -181 19 -175 53
rect -141 19 -135 53
rect -181 -19 -135 19
rect -181 -53 -175 -19
rect -141 -53 -135 -19
rect -181 -100 -135 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 135 53 181 100
rect 135 19 141 53
rect 175 19 181 53
rect 135 -19 181 19
rect 135 -53 141 -19
rect 175 -53 181 -19
rect 135 -100 181 -53
rect 293 53 339 100
rect 293 19 299 53
rect 333 19 339 53
rect 293 -19 339 19
rect 293 -53 299 -19
rect 333 -53 339 -19
rect 293 -100 339 -53
rect -283 -138 -191 -132
rect -283 -172 -254 -138
rect -220 -172 -191 -138
rect -283 -178 -191 -172
rect -125 -138 -33 -132
rect -125 -172 -96 -138
rect -62 -172 -33 -138
rect -125 -178 -33 -172
rect 33 -138 125 -132
rect 33 -172 62 -138
rect 96 -172 125 -138
rect 33 -178 125 -172
rect 191 -138 283 -132
rect 191 -172 220 -138
rect 254 -172 283 -138
rect 191 -178 283 -172
<< properties >>
string FIXED_BBOX -450 -293 450 293
<< end >>
