magic
tech sky130A
magscale 1 2
timestamp 1699617814
<< checkpaint >>
rect -1260 -1260 70034 104785
<< metal1 >>
rect 788 90615 1322 90641
rect 788 90583 801 90615
rect 784 90499 801 90583
rect 1301 90583 1322 90615
rect 1301 90499 2290 90583
rect 784 90479 2290 90499
rect 1806 87773 2212 87798
rect 1806 87529 1823 87773
rect 2195 87529 2212 87773
rect 1806 87504 2212 87529
rect 11 86970 1368 86975
rect 11 86948 1374 86970
rect 11 86832 37 86948
rect 601 86832 1374 86948
rect 11 86773 1374 86832
rect 1174 86770 1374 86773
rect 1420 84292 1702 84316
rect 1420 84048 1439 84292
rect 1683 84048 1702 84292
rect 1420 84024 1702 84048
rect 3016 83832 3316 83878
rect 3016 83204 3048 83832
rect 3292 83204 3316 83832
rect 3016 83144 3316 83204
rect 790 83005 1374 83050
rect 790 82889 825 83005
rect 1325 82889 1374 83005
rect 790 82852 1374 82889
rect 812 82850 1374 82852
rect 34580 82729 35070 82737
rect 1168 82705 1374 82714
rect 806 82671 1450 82705
rect 806 82555 844 82671
rect 1408 82555 1450 82671
rect 33304 82691 35070 82729
rect 21068 82637 21262 82641
rect 806 82521 1450 82555
rect 20506 82598 21262 82637
rect 1168 82504 1374 82521
rect 20506 82482 21109 82598
rect 21225 82482 21262 82598
rect 20506 82439 21262 82482
rect 20510 82438 20642 82439
rect 33304 82383 34639 82691
rect 35011 82383 35070 82691
rect 33304 82321 35070 82383
<< via1 >>
rect 801 90499 1301 90615
rect 1823 87529 2195 87773
rect 37 86832 601 86948
rect 1439 84048 1683 84292
rect 3048 83204 3292 83832
rect 825 82889 1325 83005
rect 844 82555 1408 82671
rect 21109 82482 21225 82598
rect 34639 82383 35011 82691
<< metal2 >>
rect 4424 103227 4520 103525
rect 7828 103225 7918 103525
rect 11230 103217 11320 103525
rect 14528 103217 14618 103525
rect 17840 103219 17936 103525
rect 21214 103219 21310 103525
rect 24516 103219 24612 103525
rect 27962 103217 28050 103525
rect 35196 103471 35256 103525
rect 35342 103471 35402 103525
rect 35488 103473 35548 103525
rect 35188 103433 35268 103471
rect 35188 103377 35203 103433
rect 35259 103377 35268 103433
rect 35188 103337 35268 103377
rect 35336 103437 35412 103471
rect 35336 103381 35346 103437
rect 35402 103381 35412 103437
rect 35336 103337 35412 103381
rect 35480 103435 35556 103473
rect 35480 103379 35494 103435
rect 35550 103379 35556 103435
rect 35480 103337 35556 103379
rect 36404 103351 36598 103525
rect 36404 103135 36426 103351
rect 36562 103135 36598 103351
rect 36404 103085 36598 103135
rect 27882 99251 28140 99307
rect 27882 99033 27899 99251
rect 27870 98795 27899 99033
rect 28115 98795 28140 99251
rect 27870 98733 28140 98795
rect 27870 98535 28132 98733
rect 788 90625 1322 90641
rect 788 90615 823 90625
rect 1279 90615 1322 90625
rect 788 90499 801 90615
rect 1301 90499 1322 90615
rect 788 90489 823 90499
rect 1279 90489 1322 90499
rect 788 90479 1322 90489
rect 1786 90405 2122 90415
rect 1786 90349 1805 90405
rect 1861 90349 1885 90405
rect 1941 90349 1965 90405
rect 2021 90349 2045 90405
rect 2101 90349 2122 90405
rect 1410 90226 1720 90246
rect 1410 90170 1455 90226
rect 1511 90170 1535 90226
rect 1591 90170 1615 90226
rect 1671 90170 1720 90226
rect 1410 87818 1720 90170
rect 1408 87488 1720 87818
rect 2 86958 632 86987
rect 2 86948 51 86958
rect 587 86948 632 86958
rect 2 86832 37 86948
rect 601 86832 632 86948
rect 2 86822 51 86832
rect 587 86822 632 86832
rect 2 86785 632 86822
rect 1410 84292 1720 87488
rect 1786 88134 2122 90349
rect 27910 90231 28132 98535
rect 27910 90175 27950 90231
rect 28006 90175 28030 90231
rect 28086 90175 28132 90231
rect 27910 90154 28132 90175
rect 3012 90039 3312 90083
rect 3012 89743 3053 90039
rect 3269 89743 3312 90039
rect 1786 87820 2240 88134
rect 1786 87773 2246 87820
rect 1786 87529 1823 87773
rect 2195 87529 2246 87773
rect 1786 87470 2246 87529
rect 1410 84048 1439 84292
rect 1683 84048 1720 84292
rect 1410 84019 1720 84048
rect 3012 83878 3312 89743
rect 3012 83832 3316 83878
rect 3012 83204 3048 83832
rect 3292 83204 3316 83832
rect 3012 83170 3316 83204
rect 3016 83144 3316 83170
rect 790 83015 1374 83050
rect 790 83005 847 83015
rect 1303 83005 1374 83015
rect 790 82889 825 83005
rect 1325 82889 1374 83005
rect 790 82879 847 82889
rect 1303 82879 1374 82889
rect 790 82852 1374 82879
rect 806 82681 1450 82705
rect 806 82671 858 82681
rect 1394 82671 1450 82681
rect 806 82555 844 82671
rect 1408 82555 1450 82671
rect 34580 82691 35070 82737
rect 34580 82685 34639 82691
rect 35011 82685 35070 82691
rect 806 82545 858 82555
rect 1394 82545 1450 82555
rect 806 82521 1450 82545
rect 21068 82608 21262 82641
rect 21068 82472 21099 82608
rect 21235 82472 21262 82608
rect 21068 82441 21262 82472
rect 34580 82389 34637 82685
rect 35013 82389 35070 82685
rect 34580 82383 34639 82389
rect 35011 82383 35070 82389
rect 34580 82329 35070 82383
rect 33630 80176 33806 80305
rect 33630 80040 33647 80176
rect 33783 80040 33806 80176
rect 33630 80009 33806 80040
rect 19202 77228 19814 77313
rect 19202 76772 19305 77228
rect 19681 76772 19814 77228
rect 19202 76703 19814 76772
rect 19346 75779 19610 76703
rect 23594 76271 24210 76339
rect 23594 75815 23659 76271
rect 24115 75815 24210 76271
rect 32200 75985 32752 75987
rect 19374 75451 19596 75779
rect 23594 75745 24210 75815
rect 32198 75896 32762 75985
rect 23770 75459 23986 75745
rect 32198 75520 32252 75896
rect 32708 75520 32762 75896
rect 32198 75447 32762 75520
rect 32200 75429 32752 75447
rect 32336 75329 32558 75429
<< via2 >>
rect 35203 103377 35259 103433
rect 35346 103381 35402 103437
rect 35494 103379 35550 103435
rect 36426 103135 36562 103351
rect 27899 98795 28115 99251
rect 823 90615 1279 90625
rect 823 90499 1279 90615
rect 823 90489 1279 90499
rect 1805 90349 1861 90405
rect 1885 90349 1941 90405
rect 1965 90349 2021 90405
rect 2045 90349 2101 90405
rect 1455 90170 1511 90226
rect 1535 90170 1591 90226
rect 1615 90170 1671 90226
rect 51 86948 587 86958
rect 51 86832 587 86948
rect 51 86822 587 86832
rect 27950 90175 28006 90231
rect 28030 90175 28086 90231
rect 3053 89743 3269 90039
rect 847 83005 1303 83015
rect 847 82889 1303 83005
rect 847 82879 1303 82889
rect 858 82671 1394 82681
rect 858 82555 1394 82671
rect 858 82545 1394 82555
rect 21099 82598 21235 82608
rect 21099 82482 21109 82598
rect 21109 82482 21225 82598
rect 21225 82482 21235 82598
rect 21099 82472 21235 82482
rect 34637 82389 34639 82685
rect 34639 82389 35011 82685
rect 35011 82389 35013 82685
rect 33647 80040 33783 80176
rect 19305 76772 19681 77228
rect 23659 75815 24115 76271
rect 32252 75520 32708 75896
<< metal3 >>
rect 35341 103471 35402 103495
rect 35488 103473 35548 103495
rect 35188 103433 35268 103471
rect 35188 103377 35203 103433
rect 35259 103377 35268 103433
rect 35188 103337 35268 103377
rect 35336 103437 35412 103471
rect 35336 103381 35346 103437
rect 35402 103381 35412 103437
rect 35336 103337 35412 103381
rect 35480 103435 35556 103473
rect 35480 103379 35494 103435
rect 35550 103379 35556 103435
rect 35480 103337 35556 103379
rect 36406 103351 36598 103405
rect 27882 99255 28140 99307
rect 27882 98791 27895 99255
rect 28119 98791 28140 99255
rect 27882 98733 28140 98791
rect 35196 97395 35256 103337
rect 34802 97335 35256 97395
rect 35341 97257 35402 103337
rect 34910 97197 35402 97257
rect 35107 97196 35402 97197
rect 35107 97195 35363 97196
rect 35488 97123 35548 103337
rect 34812 97063 35548 97123
rect 36406 103135 36426 103351
rect 36562 103135 36598 103351
rect 21304 94797 21512 94837
rect 21304 94733 21335 94797
rect 21399 94733 21415 94797
rect 21479 94733 21512 94797
rect 21304 94685 21512 94733
rect 788 90625 1322 90641
rect 788 90589 823 90625
rect 1279 90589 1322 90625
rect 788 90525 819 90589
rect 1283 90525 1322 90589
rect 788 90489 823 90525
rect 1279 90489 1322 90525
rect 788 90479 1322 90489
rect 1210 90405 36296 90417
rect 1210 90349 1805 90405
rect 1861 90349 1885 90405
rect 1941 90349 1965 90405
rect 2021 90349 2045 90405
rect 2101 90403 36296 90405
rect 2101 90349 24658 90403
rect 1210 90339 24658 90349
rect 24722 90339 24738 90403
rect 24802 90339 24818 90403
rect 24882 90339 24898 90403
rect 24962 90401 36296 90403
rect 24962 90339 34060 90401
rect 1210 90337 34060 90339
rect 34124 90337 34140 90401
rect 34204 90337 34220 90401
rect 34284 90337 34300 90401
rect 34364 90337 36296 90401
rect 1210 90323 36296 90337
rect 1206 90239 36296 90247
rect 1204 90234 36296 90239
rect 1204 90231 34594 90234
rect 1204 90226 27950 90231
rect 1204 90170 1455 90226
rect 1511 90170 1535 90226
rect 1591 90170 1615 90226
rect 1671 90175 27950 90226
rect 28006 90175 28030 90231
rect 28086 90175 34594 90231
rect 1671 90170 34594 90175
rect 34658 90170 34674 90234
rect 34738 90170 34754 90234
rect 34818 90170 34834 90234
rect 34898 90170 34914 90234
rect 34978 90170 34994 90234
rect 35058 90170 36296 90234
rect 1204 90153 36296 90170
rect 1204 90149 1502 90153
rect 1204 90083 2354 90085
rect 1200 90055 36296 90083
rect 1200 90039 35247 90055
rect 1200 89743 3053 90039
rect 3269 90038 35247 90039
rect 3269 89894 21333 90038
rect 21477 89894 35247 90038
rect 3269 89751 35247 89894
rect 35631 89751 36296 90055
rect 3269 89743 36296 89751
rect 1200 89683 36296 89743
rect 1210 89561 36296 89601
rect 1210 89291 2269 89561
rect 1224 89257 2269 89291
rect 2573 89553 36296 89561
rect 2573 89257 32676 89553
rect 1224 89249 32676 89257
rect 32820 89546 36296 89553
rect 32820 89249 35845 89546
rect 1224 89242 35845 89249
rect 36229 89242 36296 89546
rect 1224 89201 36296 89242
rect 0 86958 640 86975
rect 0 86822 51 86958
rect 587 86822 640 86958
rect 0 86773 640 86822
rect 33610 83267 34422 83323
rect 790 83019 1374 83050
rect 790 82875 843 83019
rect 1307 82875 1374 83019
rect 790 82852 1374 82875
rect 33610 82883 34064 83267
rect 34368 82883 34422 83267
rect 33610 82819 34422 82883
rect 0 82707 560 82713
rect 0 82705 1446 82707
rect 0 82685 1450 82705
rect 0 82541 854 82685
rect 1398 82541 1450 82685
rect 34580 82689 35070 82737
rect 0 82527 1450 82541
rect 806 82521 1450 82527
rect 21068 82608 21260 82657
rect 21068 82472 21099 82608
rect 21235 82472 21260 82608
rect 21068 80945 21260 82472
rect 34580 82385 34633 82689
rect 35017 82385 35070 82689
rect 34580 82329 35070 82385
rect 34798 82223 35212 82227
rect 36406 82223 36598 103135
rect 33004 82031 36598 82223
rect 34798 82029 35212 82031
rect 19202 77228 19814 77313
rect 19202 76772 19305 77228
rect 19681 77111 19814 77228
rect 21070 77111 21262 80844
rect 33630 80276 33806 80305
rect 33630 80052 33643 80276
rect 33787 80052 33806 80276
rect 33630 80040 33647 80052
rect 33783 80040 33806 80052
rect 33630 80009 33806 80040
rect 19681 76919 21262 77111
rect 19681 76772 19814 76919
rect 19202 76703 19814 76772
rect 23594 76327 24210 76339
rect 802 76323 33490 76327
rect 802 76294 33840 76323
rect 802 76150 854 76294
rect 1158 76271 33840 76294
rect 1158 76150 23659 76271
rect 802 76131 23659 76150
rect 806 76127 23659 76131
rect 23594 75815 23659 76127
rect 24115 76252 33840 76271
rect 24115 76188 33448 76252
rect 33512 76188 33528 76252
rect 33592 76188 33608 76252
rect 33672 76188 33688 76252
rect 33752 76188 33768 76252
rect 33832 76188 33840 76252
rect 24115 76127 33840 76188
rect 24115 75815 24210 76127
rect 33410 76113 33840 76127
rect 32200 75985 32752 75987
rect 23594 75745 24210 75815
rect 32198 75896 32762 75985
rect 0 75625 1624 75635
rect 32198 75625 32252 75896
rect 0 75520 32252 75625
rect 32708 75520 32762 75896
rect 0 75447 32762 75520
rect 0 75433 32752 75447
rect 32200 75429 32752 75433
rect 34048 75223 34374 75243
rect 34048 74759 34059 75223
rect 34363 74759 34374 75223
rect 34048 74739 34374 74759
rect 34598 74440 35030 74441
rect 34598 73976 34622 74440
rect 35006 73976 35030 74440
rect 34598 73975 35030 73976
rect 35258 73618 35664 73623
rect 35258 73154 35269 73618
rect 35653 73154 35664 73618
rect 35258 73149 35664 73154
rect 35826 72815 36246 72843
rect 35826 72351 35844 72815
rect 36228 72351 36246 72815
rect 35826 72323 36246 72351
rect 0 63923 2356 64099
rect 0 57197 2360 57373
rect 0 50481 2352 50657
rect 0 43787 2364 43963
rect 0 37017 2368 37193
rect 0 36105 2356 36281
rect 0 35639 2346 35815
rect 0 30031 2356 30207
rect 0 23325 2364 23501
rect 0 16605 2360 16781
rect 0 9903 2352 10079
rect 0 3125 2356 3301
rect 0 1982 888 1987
rect 1212 1982 2650 1983
rect 0 1587 2650 1982
rect 1212 1585 2650 1587
rect 0 1449 888 1451
rect 0 1051 2644 1449
rect 0 947 924 951
rect 0 559 2688 947
rect 0 376 2686 387
rect 0 0 3272 376
<< via3 >>
rect 27895 99251 28119 99255
rect 27895 98795 27899 99251
rect 27899 98795 28115 99251
rect 28115 98795 28119 99251
rect 27895 98791 28119 98795
rect 21335 94733 21399 94797
rect 21415 94733 21479 94797
rect 819 90525 823 90589
rect 823 90525 883 90589
rect 899 90525 963 90589
rect 979 90525 1043 90589
rect 1059 90525 1123 90589
rect 1139 90525 1203 90589
rect 1219 90525 1279 90589
rect 1279 90525 1283 90589
rect 24658 90339 24722 90403
rect 24738 90339 24802 90403
rect 24818 90339 24882 90403
rect 24898 90339 24962 90403
rect 34060 90337 34124 90401
rect 34140 90337 34204 90401
rect 34220 90337 34284 90401
rect 34300 90337 34364 90401
rect 34594 90170 34658 90234
rect 34674 90170 34738 90234
rect 34754 90170 34818 90234
rect 34834 90170 34898 90234
rect 34914 90170 34978 90234
rect 34994 90170 35058 90234
rect 21333 89894 21477 90038
rect 35247 89751 35631 90055
rect 2269 89257 2573 89561
rect 32676 89249 32820 89553
rect 35845 89242 36229 89546
rect 843 83015 1307 83019
rect 843 82879 847 83015
rect 847 82879 1303 83015
rect 1303 82879 1307 83015
rect 843 82875 1307 82879
rect 34064 82883 34368 83267
rect 854 82681 1398 82685
rect 854 82545 858 82681
rect 858 82545 1394 82681
rect 1394 82545 1398 82681
rect 854 82541 1398 82545
rect 34633 82685 35017 82689
rect 34633 82389 34637 82685
rect 34637 82389 35013 82685
rect 35013 82389 35017 82685
rect 34633 82385 35017 82389
rect 33643 80176 33787 80276
rect 33643 80052 33647 80176
rect 33647 80052 33783 80176
rect 33783 80052 33787 80176
rect 854 76150 1158 76294
rect 33448 76188 33512 76252
rect 33528 76188 33592 76252
rect 33608 76188 33672 76252
rect 33688 76188 33752 76252
rect 33768 76188 33832 76252
rect 34059 74759 34363 75223
rect 34622 73976 35006 74440
rect 35269 73154 35653 73618
rect 35844 72351 36228 72815
<< metal4 >>
rect 27894 99255 28120 99289
rect 27894 98791 27895 99255
rect 28119 98791 28120 99255
rect 27894 98757 28120 98791
rect 21304 94797 21512 94837
rect 21304 94733 21335 94797
rect 21399 94733 21415 94797
rect 21479 94733 21512 94797
rect 21304 94685 21512 94733
rect 788 90589 1322 90641
rect 788 90525 819 90589
rect 883 90525 899 90589
rect 963 90525 979 90589
rect 1043 90525 1059 90589
rect 1123 90525 1139 90589
rect 1203 90525 1219 90589
rect 1283 90525 1322 90589
rect 788 90479 1322 90525
rect 792 83810 992 90479
rect 21304 90038 21510 94685
rect 24650 90403 24970 98499
rect 24650 90339 24658 90403
rect 24722 90339 24738 90403
rect 24802 90339 24818 90403
rect 24882 90339 24898 90403
rect 24962 90339 24970 90403
rect 24650 90325 24970 90339
rect 34016 90401 34412 90415
rect 34016 90337 34060 90401
rect 34124 90337 34140 90401
rect 34204 90337 34220 90401
rect 34284 90337 34300 90401
rect 34364 90337 34412 90401
rect 21304 89894 21333 90038
rect 21477 89894 21510 90038
rect 2202 89561 2626 89601
rect 2202 89257 2269 89561
rect 2573 89257 2626 89561
rect 2202 88906 2626 89257
rect 2202 88633 2628 88906
rect 2208 88276 2628 88633
rect 21304 87704 21510 89894
rect 32627 89553 32861 89600
rect 32627 89249 32676 89553
rect 32820 89249 32861 89553
rect 32627 87684 32861 89249
rect 776 83384 992 83810
rect 792 83050 992 83384
rect 34016 83339 34412 90337
rect 34588 90234 35066 90424
rect 34588 90170 34594 90234
rect 34658 90170 34674 90234
rect 34738 90170 34754 90234
rect 34818 90170 34834 90234
rect 34898 90170 34914 90234
rect 34978 90170 34994 90234
rect 35058 90170 35066 90234
rect 34016 83267 34428 83339
rect 790 83019 1374 83050
rect 790 82875 843 83019
rect 1307 82875 1374 83019
rect 790 82852 1374 82875
rect 34016 82883 34064 83267
rect 34368 82883 34428 83267
rect 792 82850 1372 82852
rect 792 82848 992 82850
rect 34016 82807 34428 82883
rect 804 82705 1012 82711
rect 804 82685 1450 82705
rect 804 82541 854 82685
rect 1398 82541 1450 82685
rect 804 82521 1450 82541
rect 804 76327 1012 82521
rect 33630 80276 33810 80307
rect 33630 80052 33643 80276
rect 33787 80052 33810 80276
rect 33630 80009 33810 80052
rect 802 76294 1216 76327
rect 33630 76323 33808 80009
rect 802 76150 854 76294
rect 1158 76150 1216 76294
rect 802 76131 1216 76150
rect 33410 76252 33840 76323
rect 33410 76188 33448 76252
rect 33512 76188 33528 76252
rect 33592 76188 33608 76252
rect 33672 76188 33688 76252
rect 33752 76188 33768 76252
rect 33832 76188 33840 76252
rect 33410 76113 33840 76188
rect 34016 75223 34412 82807
rect 34016 74759 34059 75223
rect 34363 74759 34412 75223
rect 34016 74673 34412 74759
rect 34588 82741 35066 90170
rect 35204 90055 35682 90416
rect 35204 89751 35247 90055
rect 35631 89751 35682 90055
rect 34588 82689 35070 82741
rect 34588 82385 34633 82689
rect 35017 82385 35070 82689
rect 34588 82329 35070 82385
rect 34588 74440 35066 82329
rect 34588 73976 34622 74440
rect 35006 73976 35066 74440
rect 34588 73902 35066 73976
rect 35204 73618 35682 89751
rect 35204 73154 35269 73618
rect 35653 73154 35682 73618
rect 35204 73104 35682 73154
rect 35806 89546 36284 90419
rect 35806 89242 35845 89546
rect 36229 89242 36284 89546
rect 35806 72815 36284 89242
rect 35806 72351 35844 72815
rect 36228 72351 36284 72815
rect 35806 72302 36284 72351
use EF_AMUX0801WISO  EF_AMUX0801WISO_0
timestamp 1699616113
transform 1 0 1516 0 -1 101519
box -306 -2006 33704 11044
use EF_DACSCA1001  EF_DACSCA1001_0
timestamp 1699616113
transform 1 0 2156 0 1 7090
box -946 -7090 66618 68998
use EF_R2RVCE  EF_R2RVCE_0
timestamp 1699616113
transform 1 0 21872 0 1 77914
box -804 -1465 11921 11144
use sample_and_hold  sample_and_hold_0
timestamp 1699616113
transform 1 0 1174 0 1 77864
box 0 -114 19469 11183
<< labels >>
flabel metal3 s 0 86773 640 86975 0 FreeSans 235 0 0 0 HOLD
port 1 nsew
flabel metal1 s 1174 86770 1374 86970 0 FreeSans 13 0 0 0 HOLD
port 1 nsew
flabel metal2 s 27962 103217 28050 103525 0 FreeSans 60 0 0 0 VIN[0]
port 2 nsew
flabel metal2 s 24516 103219 24612 103525 0 FreeSans 60 0 0 0 VIN[1]
port 3 nsew
flabel metal2 s 21214 103219 21310 103525 0 FreeSans 60 0 0 0 VIN[2]
port 4 nsew
flabel metal2 s 17840 103219 17936 103525 0 FreeSans 60 0 0 0 VIN[3]
port 5 nsew
flabel metal2 s 14528 103217 14618 103525 0 FreeSans 60 0 0 0 VIN[4]
port 6 nsew
flabel metal2 s 11230 103217 11320 103525 0 FreeSans 60 0 0 0 VIN[5]
port 7 nsew
flabel metal2 s 7828 103225 7918 103525 0 FreeSans 60 0 0 0 VIN[6]
port 8 nsew
flabel metal2 s 4424 103227 4520 103525 0 FreeSans 60 0 0 0 VIN[7]
port 9 nsew
flabel metal3 s 0 82527 560 82713 0 FreeSans 235 0 0 0 EN
port 10 nsew
flabel metal3 s 0 75433 500 75635 0 FreeSans 235 0 0 0 RST
port 11 nsew
flabel metal3 s 0 63923 554 64099 0 FreeSans 235 0 0 0 DATA[9]
port 12 nsew
flabel metal3 s 0 57197 648 57373 0 FreeSans 235 0 0 0 DATA[8]
port 13 nsew
flabel metal3 s 0 50481 648 50657 0 FreeSans 235 0 0 0 DATA[7]
port 14 nsew
flabel metal3 s 0 43787 648 43963 0 FreeSans 235 0 0 0 DATA[6]
port 15 nsew
flabel metal3 s 0 37017 648 37193 0 FreeSans 235 0 0 0 DATA[5]
port 16 nsew
flabel metal3 s 0 30031 648 30207 0 FreeSans 235 0 0 0 DATA[0]
port 17 nsew
flabel metal3 s 0 23325 648 23501 0 FreeSans 235 0 0 0 DATA[1]
port 18 nsew
flabel metal3 s 0 16605 648 16781 0 FreeSans 235 0 0 0 DATA[2]
port 19 nsew
flabel metal3 s 0 9903 648 10079 0 FreeSans 235 0 0 0 DATA[3]
port 20 nsew
flabel metal3 s 0 3125 648 3301 0 FreeSans 235 0 0 0 DATA[4]
port 21 nsew
flabel metal3 s 0 1051 888 1451 0 FreeSans 235 0 0 0 DVSS
port 22 nsew
flabel metal3 s 0 1587 888 1987 0 FreeSans 235 0 0 0 DVDD
port 23 nsew
flabel metal3 s 0 559 924 951 0 FreeSans 235 0 0 0 VDD
port 24 nsew
flabel metal3 s 0 36105 658 36281 0 FreeSans 235 0 0 0 VH
port 25 nsew
flabel metal3 s 0 35639 658 35815 0 FreeSans 235 0 0 0 VL
port 26 nsew
flabel metal2 s 35196 103341 35256 103525 0 FreeSans 235 0 0 0 B[0]
port 27 nsew
flabel metal2 s 35342 103337 35402 103525 0 FreeSans 235 0 0 0 B[1]
port 28 nsew
flabel metal2 s 35488 103337 35548 103525 0 FreeSans 235 0 0 0 B[2]
port 29 nsew
flabel metal2 s 36404 103085 36598 103525 0 FreeSans 235 0 0 0 CMP
port 30 nsew
flabel metal3 s 0 0 1224 386 0 FreeSans 600 0 0 0 VSS
port 31 nsew
<< end >>
