VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO EF_ADCS1008NC
  CLASS BLOCK ;
  FOREIGN EF_ADCS1008NC ;
  ORIGIN 0.000 0.000 ;
  SIZE 343.870 BY 518.865 ;
  PIN HOLD
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT 5.870 435.090 6.870 436.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 435.105 3.200 436.115 ;
    END
  END HOLD
  PIN VIN[0]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 139.810 517.325 140.250 518.865 ;
    END
  END VIN[0]
  PIN VIN[1]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 122.580 517.335 123.060 518.865 ;
    END
  END VIN[1]
  PIN VIN[2]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 106.070 517.335 106.550 518.865 ;
    END
  END VIN[2]
  PIN VIN[3]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 89.200 517.335 89.680 518.865 ;
    END
  END VIN[3]
  PIN VIN[4]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 72.640 517.325 73.090 518.865 ;
    END
  END VIN[4]
  PIN VIN[5]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 56.150 517.325 56.600 518.865 ;
    END
  END VIN[5]
  PIN VIN[6]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 39.140 517.365 39.590 518.865 ;
    END
  END VIN[6]
  PIN VIN[7]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 22.120 517.375 22.600 518.865 ;
    END
  END VIN[7]
  PIN EN
    ANTENNAGATEAREA 1.752000 ;
    ANTENNADIFFAREA 1.080000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.875 2.800 414.805 ;
    END
  END EN
  PIN RST
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.405 2.500 379.415 ;
    END
  END RST
  PIN DATA[9]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.855 2.770 321.735 ;
    END
  END DATA[9]
  PIN DATA[8]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.225 3.240 288.105 ;
    END
  END DATA[8]
  PIN DATA[7]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.645 3.240 254.525 ;
    END
  END DATA[7]
  PIN DATA[6]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.175 3.240 221.055 ;
    END
  END DATA[6]
  PIN DATA[5]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.325 3.240 187.205 ;
    END
  END DATA[5]
  PIN DATA[0]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.395 3.240 152.275 ;
    END
  END DATA[0]
  PIN DATA[1]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.865 3.240 118.745 ;
    END
  END DATA[1]
  PIN DATA[2]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.265 3.240 85.145 ;
    END
  END DATA[2]
  PIN DATA[3]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.755 3.240 51.635 ;
    END
  END DATA[3]
  PIN DATA[4]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.865 3.240 17.745 ;
    END
  END DATA[4]
  PIN DVSS
    ANTENNAGATEAREA 74.759102 ;
    ANTENNADIFFAREA 1023.766663 ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.495 4.440 8.495 ;
    END
  END DVSS
  PIN DVDD
    ANTENNAGATEAREA 47.261497 ;
    ANTENNADIFFAREA 93.596451 ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.175 4.440 11.175 ;
    END
  END DVDD
  PIN VDD
    ANTENNAGATEAREA 100.000000 ;
    ANTENNADIFFAREA 2509.495605 ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.035 4.620 5.995 ;
    END
  END VDD
  PIN VSS
    ANTENNAGATEAREA 130.500000 ;
    ANTENNADIFFAREA 621.362671 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.275 4.700 3.175 ;
    END
  END VSS
  PIN VH
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.765 3.290 182.645 ;
    END
  END VH
  PIN VL
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.435 3.290 180.315 ;
    END
  END VL
  PIN B[0]
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 175.980 517.945 176.280 518.865 ;
    END
  END B[0]
  PIN B[1]
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 176.710 517.925 177.010 518.865 ;
    END
  END B[1]
  PIN B[2]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 177.440 517.925 177.740 518.865 ;
    END
  END B[2]
  PIN CMP
    ANTENNADIFFAREA 0.492900 ;
    PORT
      LAYER met2 ;
        RECT 182.020 516.665 182.990 518.865 ;
    END
  END CMP
  OBS
      LAYER li1 ;
        RECT 7.235 15.315 247.920 508.630 ;
      LAYER met1 ;
        RECT 0.055 436.370 248.615 508.835 ;
        RECT 0.055 434.810 5.590 436.370 ;
        RECT 7.150 434.810 248.615 436.370 ;
        RECT 0.055 13.000 248.615 434.810 ;
      LAYER met2 ;
        RECT 0.010 517.095 21.840 518.840 ;
        RECT 22.880 517.095 38.860 518.840 ;
        RECT 0.010 517.085 38.860 517.095 ;
        RECT 39.870 517.085 55.870 518.840 ;
        RECT 0.010 517.045 55.870 517.085 ;
        RECT 56.880 517.045 72.360 518.840 ;
        RECT 73.370 517.055 88.920 518.840 ;
        RECT 89.960 517.055 105.790 518.840 ;
        RECT 106.830 517.055 122.300 518.840 ;
        RECT 123.340 517.055 139.530 518.840 ;
        RECT 73.370 517.045 139.530 517.055 ;
        RECT 140.530 517.665 175.700 518.840 ;
        RECT 140.530 517.645 176.430 517.665 ;
        RECT 178.020 517.645 181.740 518.840 ;
        RECT 140.530 517.045 181.740 517.645 ;
        RECT 0.010 516.385 181.740 517.045 ;
        RECT 183.270 516.385 246.300 518.840 ;
        RECT 0.010 13.000 246.300 516.385 ;
      LAYER met3 ;
        RECT 2.500 436.515 343.870 518.715 ;
        RECT 3.600 434.705 343.870 436.515 ;
        RECT 2.500 415.205 343.870 434.705 ;
        RECT 3.200 413.475 343.870 415.205 ;
        RECT 2.500 379.815 343.870 413.475 ;
        RECT 2.900 378.005 343.870 379.815 ;
        RECT 2.500 322.135 343.870 378.005 ;
        RECT 3.170 320.455 343.870 322.135 ;
        RECT 2.500 288.505 343.870 320.455 ;
        RECT 3.640 286.825 343.870 288.505 ;
        RECT 2.500 254.925 343.870 286.825 ;
        RECT 3.640 253.245 343.870 254.925 ;
        RECT 2.500 221.455 343.870 253.245 ;
        RECT 3.640 219.775 343.870 221.455 ;
        RECT 2.500 187.605 343.870 219.775 ;
        RECT 3.640 185.925 343.870 187.605 ;
        RECT 2.500 183.045 343.870 185.925 ;
        RECT 3.690 181.365 343.870 183.045 ;
        RECT 2.500 180.715 343.870 181.365 ;
        RECT 3.690 179.035 343.870 180.715 ;
        RECT 2.500 152.675 343.870 179.035 ;
        RECT 3.640 150.995 343.870 152.675 ;
        RECT 2.500 119.145 343.870 150.995 ;
        RECT 3.640 117.465 343.870 119.145 ;
        RECT 2.500 85.545 343.870 117.465 ;
        RECT 3.640 83.865 343.870 85.545 ;
        RECT 2.500 52.035 343.870 83.865 ;
        RECT 3.640 50.355 343.870 52.035 ;
        RECT 2.500 18.145 343.870 50.355 ;
        RECT 3.640 16.465 343.870 18.145 ;
        RECT 2.500 11.575 343.870 16.465 ;
        RECT 4.840 6.395 343.870 11.575 ;
        RECT 5.020 3.635 343.870 6.395 ;
        RECT 2.500 3.575 343.870 3.635 ;
        RECT 5.100 1.240 343.870 3.575 ;
      LAYER met4 ;
        RECT 3.880 1.240 343.700 516.835 ;
      LAYER met5 ;
        RECT 16.945 385.720 170.975 508.150 ;
  END
END EF_ADCS1008NC
END LIBRARY

