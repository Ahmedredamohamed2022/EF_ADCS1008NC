magic
tech sky130A
timestamp 1699926577
use sky130_fd_pr__cap_mim_m3_1_STW68H  sky130_fd_pr__cap_mim_m3_1_STW68H_0
timestamp 1699926577
transform -1 0 1243 0 1 520
box -1243 -520 1243 520
use sky130_fd_pr__cap_mim_m3_1_STW68H  sky130_fd_pr__cap_mim_m3_1_STW68H_1
timestamp 1699926577
transform -1 0 4243 0 1 520
box -1243 -520 1243 520
use sky130_fd_pr__cap_mim_m3_1_STW68H  sky130_fd_pr__cap_mim_m3_1_STW68H_2
timestamp 1699926577
transform -1 0 7243 0 1 520
box -1243 -520 1243 520
use sky130_fd_pr__cap_mim_m3_1_STW68H  sky130_fd_pr__cap_mim_m3_1_STW68H_3
timestamp 1699926577
transform -1 0 10243 0 1 520
box -1243 -520 1243 520
use sky130_fd_pr__cap_mim_m3_1_STW68H  sky130_fd_pr__cap_mim_m3_1_STW68H_4
timestamp 1699926577
transform -1 0 13243 0 1 520
box -1243 -520 1243 520
use sky130_fd_pr__cap_mim_m3_1_STW68H  sky130_fd_pr__cap_mim_m3_1_STW68H_5
timestamp 1699926577
transform -1 0 16243 0 1 520
box -1243 -520 1243 520
use sky130_fd_pr__cap_mim_m3_1_STW68H  sky130_fd_pr__cap_mim_m3_1_STW68H_6
timestamp 1699926577
transform -1 0 19243 0 1 520
box -1243 -520 1243 520
use sky130_fd_pr__cap_mim_m3_1_STW68H  sky130_fd_pr__cap_mim_m3_1_STW68H_7
timestamp 1699926577
transform -1 0 22243 0 1 520
box -1243 -520 1243 520
<< end >>
