magic
tech sky130A
magscale 1 2
timestamp 1693827120
<< metal1 >>
rect 3532 6232 7054 6424
rect 3532 6000 3724 6232
rect 6862 5790 7054 6232
rect 5980 2756 6176 3092
rect 9322 2768 9512 3396
rect 3728 686 3946 734
rect 3728 570 3766 686
rect 3882 570 3946 686
rect 3728 530 3946 570
rect 7074 713 7292 760
rect 7074 597 7123 713
rect 7239 597 7292 713
rect 7074 552 7292 597
rect 5470 205 7094 409
rect 6340 128 7002 154
rect 6340 12 6394 128
rect 6958 12 7002 128
rect 6340 6 7002 12
rect 6370 -2 6988 6
rect 3732 -198 3906 -166
rect 3732 -362 3762 -198
rect 3370 -442 3762 -362
rect 3878 -362 3906 -198
rect 3878 -442 6424 -362
rect 7086 -376 7272 -374
rect 6932 -378 7272 -376
rect 6932 -430 7120 -378
rect 7172 -430 7184 -378
rect 7236 -430 7272 -378
rect 6932 -436 7272 -430
rect 7086 -438 7272 -436
rect 3370 -476 6424 -442
rect 3370 -480 4138 -476
rect 9294 -626 9540 486
rect 6786 -790 9546 -626
<< via1 >>
rect 3766 570 3882 686
rect 7123 597 7239 713
rect 6394 12 6958 128
rect 3762 -442 3878 -198
rect 7120 -430 7172 -378
rect 7184 -430 7236 -378
<< metal2 >>
rect 7132 760 7260 766
rect 3728 686 3946 734
rect 3728 570 3766 686
rect 3882 570 3946 686
rect 3728 530 3946 570
rect 7074 713 7292 760
rect 7074 597 7123 713
rect 7239 597 7292 713
rect 7074 552 7292 597
rect 3738 -198 3910 530
rect 6340 128 7002 154
rect 6340 12 6394 128
rect 6958 12 7002 128
rect 6340 6 7002 12
rect 6370 2 6988 6
rect 3738 -342 3762 -198
rect 3732 -442 3762 -342
rect 3878 -414 3910 -198
rect 7132 -374 7260 552
rect 7086 -378 7272 -374
rect 3878 -442 3906 -414
rect 7086 -430 7120 -378
rect 7172 -430 7184 -378
rect 7236 -430 7272 -378
rect 7086 -438 7272 -430
rect 3732 -476 3906 -442
<< via2 >>
rect 6408 42 6464 98
rect 6488 42 6544 98
rect 6568 42 6624 98
rect 6648 42 6704 98
rect 6728 42 6784 98
rect 6808 42 6864 98
rect 6888 42 6944 98
<< metal3 >>
rect 4837 4067 9993 4293
rect 6464 962 6644 964
rect 4487 804 7811 962
rect 6464 154 6644 804
rect 6340 98 7002 154
rect 6340 42 6408 98
rect 6464 42 6488 98
rect 6544 42 6568 98
rect 6624 42 6648 98
rect 6704 42 6728 98
rect 6784 42 6808 98
rect 6864 42 6888 98
rect 6944 42 7002 98
rect 6340 6 7002 42
rect 6370 2 6988 6
use array_1ls_1tgm  array_1ls_1tgm_0
timestamp 1693827120
transform 1 0 6710 0 1 226
box 0 0 3070 6017
use array_1ls_1tgm  array_1ls_1tgm_1
timestamp 1693827120
transform 1 0 3364 0 1 205
box 0 0 3070 6017
use invm  invm_0
timestamp 1693827120
transform 1 0 4208 0 1 -1100
box 2164 308 2788 1248
<< labels >>
flabel metal1 s 6000 6288 6048 6348 0 FreeSans 161 0 0 0 vo
port 1 nsew
flabel metal3 s 9452 4136 9500 4196 0 FreeSans 161 0 0 0 vdd3p3
port 2 nsew
flabel metal3 s 6586 866 6616 898 0 FreeSans 161 0 0 0 vdd1p8
port 3 nsew
flabel metal1 s 6408 250 6438 284 0 FreeSans 161 0 0 0 vss
port 4 nsew
flabel metal1 s 6054 2844 6086 2912 0 FreeSans 161 0 0 0 a
port 5 nsew
flabel metal1 s 9394 2982 9448 3062 0 FreeSans 161 0 0 0 b
port 6 nsew
flabel metal1 s 3462 -438 3528 -380 0 FreeSans 161 0 0 0 sel
port 7 nsew
<< end >>
