magic
tech sky130A
magscale 1 2
timestamp 1699926577
<< metal3 >>
rect -2460 29356 49404 29556
rect -3400 27982 50400 27998
rect -3400 27838 2283 27982
rect 2907 27978 20289 27982
rect 2907 27937 8289 27978
rect 2907 27873 5056 27937
rect 5120 27873 5136 27937
rect 5200 27873 5216 27937
rect 5280 27873 5296 27937
rect 5360 27873 5376 27937
rect 5440 27873 5456 27937
rect 5520 27873 5536 27937
rect 5600 27873 5616 27937
rect 5680 27873 5696 27937
rect 5760 27873 8289 27937
rect 2907 27838 8289 27873
rect -3400 27834 8289 27838
rect 8913 27956 20289 27978
rect 8913 27834 14301 27956
rect -3400 27812 14301 27834
rect 14925 27838 20289 27956
rect 20913 27978 38263 27982
rect 20913 27968 32321 27978
rect 20913 27838 26283 27968
rect 14925 27824 26283 27838
rect 26907 27834 32321 27968
rect 32945 27838 38263 27978
rect 38887 27974 50400 27982
rect 38887 27838 44259 27974
rect 32945 27834 44259 27838
rect 26907 27830 44259 27834
rect 44883 27830 50400 27974
rect 26907 27824 50400 27830
rect 14925 27812 50400 27824
rect -3400 27792 50400 27812
rect -3198 16828 -2386 16836
rect -3208 16772 50225 16828
rect -3208 16760 17624 16772
rect -3208 16756 5640 16760
rect -3208 16692 -348 16756
rect -284 16692 -268 16756
rect -204 16692 -188 16756
rect -124 16692 -108 16756
rect -44 16692 -28 16756
rect 36 16692 52 16756
rect 116 16692 132 16756
rect 196 16692 212 16756
rect 276 16692 292 16756
rect 356 16696 5640 16756
rect 5704 16696 5720 16760
rect 5784 16696 5800 16760
rect 5864 16696 5880 16760
rect 5944 16696 5960 16760
rect 6024 16696 6040 16760
rect 6104 16696 6120 16760
rect 6184 16696 6200 16760
rect 6264 16696 6280 16760
rect 6344 16756 17624 16760
rect 6344 16696 11628 16756
rect 356 16692 11628 16696
rect 11692 16692 11708 16756
rect 11772 16692 11788 16756
rect 11852 16692 11868 16756
rect 11932 16692 11948 16756
rect 12012 16692 12028 16756
rect 12092 16692 12108 16756
rect 12172 16692 12188 16756
rect 12252 16692 12268 16756
rect 12332 16708 17624 16756
rect 17688 16708 17704 16772
rect 17768 16708 17784 16772
rect 17848 16708 17864 16772
rect 17928 16708 17944 16772
rect 18008 16708 18024 16772
rect 18088 16708 18104 16772
rect 18168 16708 18184 16772
rect 18248 16708 18264 16772
rect 18328 16764 50225 16772
rect 18328 16756 29646 16764
rect 18328 16708 23650 16756
rect 12332 16692 23650 16708
rect 23714 16692 23730 16756
rect 23794 16692 23810 16756
rect 23874 16692 23890 16756
rect 23954 16692 23970 16756
rect 24034 16692 24050 16756
rect 24114 16692 24130 16756
rect 24194 16692 24210 16756
rect 24274 16692 24290 16756
rect 24354 16700 29646 16756
rect 29710 16700 29726 16764
rect 29790 16700 29806 16764
rect 29870 16700 29886 16764
rect 29950 16700 29966 16764
rect 30030 16700 30046 16764
rect 30110 16700 30126 16764
rect 30190 16700 30206 16764
rect 30270 16700 30286 16764
rect 30350 16760 50225 16764
rect 30350 16748 41656 16760
rect 30350 16700 35622 16748
rect 24354 16692 35622 16700
rect -3208 16684 35622 16692
rect 35686 16684 35702 16748
rect 35766 16684 35782 16748
rect 35846 16684 35862 16748
rect 35926 16684 35942 16748
rect 36006 16684 36022 16748
rect 36086 16684 36102 16748
rect 36166 16684 36182 16748
rect 36246 16684 36262 16748
rect 36326 16696 41656 16748
rect 41720 16696 41736 16760
rect 41800 16696 41816 16760
rect 41880 16696 41896 16760
rect 41960 16696 41976 16760
rect 42040 16696 42056 16760
rect 42120 16696 42136 16760
rect 42200 16696 42216 16760
rect 42280 16696 42296 16760
rect 42360 16696 50225 16760
rect 36326 16684 50225 16696
rect -3208 16626 50225 16684
rect -3198 16624 -2386 16626
rect -3192 16426 -2380 16442
rect -3194 16361 50219 16426
rect -3194 16297 -351 16361
rect -287 16297 -271 16361
rect -207 16297 -191 16361
rect -127 16297 -111 16361
rect -47 16297 -31 16361
rect 33 16297 49 16361
rect 113 16297 129 16361
rect 193 16297 209 16361
rect 273 16297 289 16361
rect 353 16353 35643 16361
rect 353 16349 11635 16353
rect 353 16297 5631 16349
rect -3194 16285 5631 16297
rect 5695 16285 5711 16349
rect 5775 16285 5791 16349
rect 5855 16285 5871 16349
rect 5935 16285 5951 16349
rect 6015 16285 6031 16349
rect 6095 16285 6111 16349
rect 6175 16285 6191 16349
rect 6255 16285 6271 16349
rect 6335 16289 11635 16349
rect 11699 16289 11715 16353
rect 11779 16289 11795 16353
rect 11859 16289 11875 16353
rect 11939 16289 11955 16353
rect 12019 16289 12035 16353
rect 12099 16289 12115 16353
rect 12179 16289 12195 16353
rect 12259 16289 12275 16353
rect 12339 16349 23657 16353
rect 12339 16289 17639 16349
rect 6335 16285 17639 16289
rect 17703 16285 17719 16349
rect 17783 16285 17799 16349
rect 17863 16285 17879 16349
rect 17943 16285 17959 16349
rect 18023 16285 18039 16349
rect 18103 16285 18119 16349
rect 18183 16285 18199 16349
rect 18263 16285 18279 16349
rect 18343 16289 23657 16349
rect 23721 16289 23737 16353
rect 23801 16289 23817 16353
rect 23881 16289 23897 16353
rect 23961 16289 23977 16353
rect 24041 16289 24057 16353
rect 24121 16289 24137 16353
rect 24201 16289 24217 16353
rect 24281 16289 24297 16353
rect 24361 16289 29637 16353
rect 29701 16289 29717 16353
rect 29781 16289 29797 16353
rect 29861 16289 29877 16353
rect 29941 16289 29957 16353
rect 30021 16289 30037 16353
rect 30101 16289 30117 16353
rect 30181 16289 30197 16353
rect 30261 16289 30277 16353
rect 30341 16297 35643 16353
rect 35707 16297 35723 16361
rect 35787 16297 35803 16361
rect 35867 16297 35883 16361
rect 35947 16297 35963 16361
rect 36027 16297 36043 16361
rect 36107 16297 36123 16361
rect 36187 16297 36203 16361
rect 36267 16297 36283 16361
rect 36347 16349 50219 16361
rect 36347 16297 41639 16349
rect 30341 16289 41639 16297
rect 18343 16285 41639 16289
rect 41703 16285 41719 16349
rect 41783 16285 41799 16349
rect 41863 16285 41879 16349
rect 41943 16285 41959 16349
rect 42023 16285 42039 16349
rect 42103 16285 42119 16349
rect 42183 16285 42199 16349
rect 42263 16285 42279 16349
rect 42343 16285 50219 16349
rect -3194 16224 50219 16285
rect -3194 11116 -2370 11130
rect -3200 11106 50194 11116
rect -3200 11102 41627 11106
rect -3200 10958 23635 11102
rect 24339 11094 41627 11102
rect 24339 10958 29629 11094
rect -3200 10950 29629 10958
rect 30333 11082 41627 11094
rect 30333 10950 35599 11082
rect -3200 10938 35599 10950
rect 36303 10962 41627 11082
rect 42331 10962 50194 11106
rect 36303 10938 50194 10962
rect -3200 10912 50194 10938
rect -3214 10722 -2390 10734
rect -3214 10694 50202 10722
rect -3214 10674 17633 10694
rect -3214 10530 11663 10674
rect 12367 10550 17633 10674
rect 18337 10550 50202 10694
rect 12367 10530 50202 10550
rect -3214 10524 50202 10530
rect -3208 10518 50202 10524
rect -3408 5402 -2552 5410
rect -3414 5368 50204 5402
rect -3414 5224 5640 5368
rect 6344 5224 50204 5368
rect -3414 5198 50204 5224
rect -3414 5002 50220 5006
rect -3422 4986 50220 5002
rect -3422 4842 5652 4986
rect 6356 4842 50220 4986
rect -3422 4806 50220 4842
rect -3414 4802 50220 4806
rect -3346 2148 114 2346
rect -3406 -202 -2580 -200
rect -3406 -261 50190 -202
rect -3406 -273 17636 -261
rect -3406 -337 11648 -273
rect 11712 -337 11728 -273
rect 11792 -337 11808 -273
rect 11872 -337 11888 -273
rect 11952 -337 11968 -273
rect 12032 -337 12048 -273
rect 12112 -337 12128 -273
rect 12192 -337 12208 -273
rect 12272 -337 12288 -273
rect 12352 -325 17636 -273
rect 17700 -325 17716 -261
rect 17780 -325 17796 -261
rect 17860 -325 17876 -261
rect 17940 -325 17956 -261
rect 18020 -325 18036 -261
rect 18100 -325 18116 -261
rect 18180 -325 18196 -261
rect 18260 -325 18276 -261
rect 18340 -325 50190 -261
rect 12352 -337 50190 -325
rect -3406 -400 50190 -337
rect -3414 -602 -2588 -596
rect -3414 -622 50190 -602
rect -3414 -766 23745 -622
rect 24449 -642 35651 -622
rect 24449 -766 29807 -642
rect -3414 -786 29807 -766
rect 30511 -766 35651 -642
rect 36355 -630 50190 -622
rect 36355 -766 41653 -630
rect 30511 -774 41653 -766
rect 42357 -774 50190 -630
rect 30511 -786 50190 -774
rect -3414 -796 50190 -786
rect -3406 -800 50190 -796
rect -3208 -5917 50202 -5868
rect -3208 -5939 5690 -5917
rect -3208 -6003 -332 -5939
rect -268 -6003 -252 -5939
rect -188 -6003 -172 -5939
rect -108 -6003 -92 -5939
rect -28 -6003 -12 -5939
rect 52 -6003 68 -5939
rect 132 -6003 148 -5939
rect 212 -6003 228 -5939
rect 292 -5981 5690 -5939
rect 5754 -5981 5770 -5917
rect 5834 -5981 5850 -5917
rect 5914 -5981 5930 -5917
rect 5994 -5981 6010 -5917
rect 6074 -5981 6090 -5917
rect 6154 -5981 6170 -5917
rect 6234 -5981 6250 -5917
rect 6314 -5921 50202 -5917
rect 6314 -5923 35686 -5921
rect 6314 -5927 29646 -5923
rect 6314 -5981 11686 -5927
rect 292 -5991 11686 -5981
rect 11750 -5991 11766 -5927
rect 11830 -5991 11846 -5927
rect 11910 -5991 11926 -5927
rect 11990 -5991 12006 -5927
rect 12070 -5991 12086 -5927
rect 12150 -5991 12166 -5927
rect 12230 -5991 12246 -5927
rect 12310 -5931 29646 -5927
rect 12310 -5991 17686 -5931
rect 292 -5995 17686 -5991
rect 17750 -5995 17766 -5931
rect 17830 -5995 17846 -5931
rect 17910 -5995 17926 -5931
rect 17990 -5995 18006 -5931
rect 18070 -5995 18086 -5931
rect 18150 -5995 18166 -5931
rect 18230 -5995 18246 -5931
rect 18310 -5995 23708 -5931
rect 23772 -5995 23788 -5931
rect 23852 -5995 23868 -5931
rect 23932 -5995 23948 -5931
rect 24012 -5995 24028 -5931
rect 24092 -5995 24108 -5931
rect 24172 -5995 24188 -5931
rect 24252 -5995 24268 -5931
rect 24332 -5987 29646 -5931
rect 29710 -5987 29726 -5923
rect 29790 -5987 29806 -5923
rect 29870 -5987 29886 -5923
rect 29950 -5987 29966 -5923
rect 30030 -5987 30046 -5923
rect 30110 -5987 30126 -5923
rect 30190 -5987 30206 -5923
rect 30270 -5985 35686 -5923
rect 35750 -5985 35766 -5921
rect 35830 -5985 35846 -5921
rect 35910 -5985 35926 -5921
rect 35990 -5985 36006 -5921
rect 36070 -5985 36086 -5921
rect 36150 -5985 36166 -5921
rect 36230 -5985 36246 -5921
rect 36310 -5939 50202 -5921
rect 36310 -5985 41652 -5939
rect 30270 -5987 41652 -5985
rect 24332 -5995 41652 -5987
rect 292 -6003 41652 -5995
rect 41716 -6003 41732 -5939
rect 41796 -6003 41812 -5939
rect 41876 -6003 41892 -5939
rect 41956 -6003 41972 -5939
rect 42036 -6003 42052 -5939
rect 42116 -6003 42132 -5939
rect 42196 -6003 42212 -5939
rect 42276 -6003 50202 -5939
rect -3208 -6068 50202 -6003
rect -3204 -6320 50186 -6312
rect -3204 -6350 5655 -6320
rect -3204 -6494 -335 -6350
rect 369 -6464 5655 -6350
rect 6359 -6464 11635 -6320
rect 12339 -6346 23647 -6320
rect 12339 -6464 17639 -6346
rect 369 -6490 17639 -6464
rect 18343 -6464 23647 -6346
rect 24351 -6324 50186 -6320
rect 24351 -6336 41643 -6324
rect 24351 -6464 29647 -6336
rect 18343 -6480 29647 -6464
rect 30351 -6340 41643 -6336
rect 30351 -6480 35631 -6340
rect 18343 -6484 35631 -6480
rect 36335 -6468 41643 -6340
rect 42347 -6468 50186 -6324
rect 36335 -6484 50186 -6468
rect 18343 -6490 50186 -6484
rect 369 -6494 50186 -6490
rect -3204 -6512 50186 -6494
rect -3399 -17444 50401 -17426
rect -3399 -17448 20255 -17444
rect -3399 -17458 14263 -17448
rect -3399 -17602 -922 -17458
rect -298 -17460 8313 -17458
rect -298 -17602 2245 -17460
rect -3399 -17604 2245 -17602
rect 2949 -17602 8313 -17460
rect 9017 -17592 14263 -17458
rect 14967 -17588 20255 -17448
rect 20959 -17446 50401 -17444
rect 20959 -17588 26225 -17446
rect 14967 -17590 26225 -17588
rect 26929 -17450 50401 -17446
rect 26929 -17456 38251 -17450
rect 26929 -17590 32245 -17456
rect 14967 -17592 32245 -17590
rect 9017 -17600 32245 -17592
rect 32949 -17594 38251 -17456
rect 38955 -17456 50401 -17450
rect 38955 -17594 44237 -17456
rect 32949 -17600 44237 -17594
rect 44941 -17600 50401 -17456
rect 9017 -17602 50401 -17600
rect 2949 -17604 50401 -17602
rect -3399 -17632 50401 -17604
rect 5142 -19000 5782 -18970
rect -2177 -19206 49383 -19000
<< via3 >>
rect 2283 27838 2907 27982
rect 5056 27873 5120 27937
rect 5136 27873 5200 27937
rect 5216 27873 5280 27937
rect 5296 27873 5360 27937
rect 5376 27873 5440 27937
rect 5456 27873 5520 27937
rect 5536 27873 5600 27937
rect 5616 27873 5680 27937
rect 5696 27873 5760 27937
rect 8289 27834 8913 27978
rect 14301 27812 14925 27956
rect 20289 27838 20913 27982
rect 26283 27824 26907 27968
rect 32321 27834 32945 27978
rect 38263 27838 38887 27982
rect 44259 27830 44883 27974
rect -348 16692 -284 16756
rect -268 16692 -204 16756
rect -188 16692 -124 16756
rect -108 16692 -44 16756
rect -28 16692 36 16756
rect 52 16692 116 16756
rect 132 16692 196 16756
rect 212 16692 276 16756
rect 292 16692 356 16756
rect 5640 16696 5704 16760
rect 5720 16696 5784 16760
rect 5800 16696 5864 16760
rect 5880 16696 5944 16760
rect 5960 16696 6024 16760
rect 6040 16696 6104 16760
rect 6120 16696 6184 16760
rect 6200 16696 6264 16760
rect 6280 16696 6344 16760
rect 11628 16692 11692 16756
rect 11708 16692 11772 16756
rect 11788 16692 11852 16756
rect 11868 16692 11932 16756
rect 11948 16692 12012 16756
rect 12028 16692 12092 16756
rect 12108 16692 12172 16756
rect 12188 16692 12252 16756
rect 12268 16692 12332 16756
rect 17624 16708 17688 16772
rect 17704 16708 17768 16772
rect 17784 16708 17848 16772
rect 17864 16708 17928 16772
rect 17944 16708 18008 16772
rect 18024 16708 18088 16772
rect 18104 16708 18168 16772
rect 18184 16708 18248 16772
rect 18264 16708 18328 16772
rect 23650 16692 23714 16756
rect 23730 16692 23794 16756
rect 23810 16692 23874 16756
rect 23890 16692 23954 16756
rect 23970 16692 24034 16756
rect 24050 16692 24114 16756
rect 24130 16692 24194 16756
rect 24210 16692 24274 16756
rect 24290 16692 24354 16756
rect 29646 16700 29710 16764
rect 29726 16700 29790 16764
rect 29806 16700 29870 16764
rect 29886 16700 29950 16764
rect 29966 16700 30030 16764
rect 30046 16700 30110 16764
rect 30126 16700 30190 16764
rect 30206 16700 30270 16764
rect 30286 16700 30350 16764
rect 35622 16684 35686 16748
rect 35702 16684 35766 16748
rect 35782 16684 35846 16748
rect 35862 16684 35926 16748
rect 35942 16684 36006 16748
rect 36022 16684 36086 16748
rect 36102 16684 36166 16748
rect 36182 16684 36246 16748
rect 36262 16684 36326 16748
rect 41656 16696 41720 16760
rect 41736 16696 41800 16760
rect 41816 16696 41880 16760
rect 41896 16696 41960 16760
rect 41976 16696 42040 16760
rect 42056 16696 42120 16760
rect 42136 16696 42200 16760
rect 42216 16696 42280 16760
rect 42296 16696 42360 16760
rect -351 16297 -287 16361
rect -271 16297 -207 16361
rect -191 16297 -127 16361
rect -111 16297 -47 16361
rect -31 16297 33 16361
rect 49 16297 113 16361
rect 129 16297 193 16361
rect 209 16297 273 16361
rect 289 16297 353 16361
rect 5631 16285 5695 16349
rect 5711 16285 5775 16349
rect 5791 16285 5855 16349
rect 5871 16285 5935 16349
rect 5951 16285 6015 16349
rect 6031 16285 6095 16349
rect 6111 16285 6175 16349
rect 6191 16285 6255 16349
rect 6271 16285 6335 16349
rect 11635 16289 11699 16353
rect 11715 16289 11779 16353
rect 11795 16289 11859 16353
rect 11875 16289 11939 16353
rect 11955 16289 12019 16353
rect 12035 16289 12099 16353
rect 12115 16289 12179 16353
rect 12195 16289 12259 16353
rect 12275 16289 12339 16353
rect 17639 16285 17703 16349
rect 17719 16285 17783 16349
rect 17799 16285 17863 16349
rect 17879 16285 17943 16349
rect 17959 16285 18023 16349
rect 18039 16285 18103 16349
rect 18119 16285 18183 16349
rect 18199 16285 18263 16349
rect 18279 16285 18343 16349
rect 23657 16289 23721 16353
rect 23737 16289 23801 16353
rect 23817 16289 23881 16353
rect 23897 16289 23961 16353
rect 23977 16289 24041 16353
rect 24057 16289 24121 16353
rect 24137 16289 24201 16353
rect 24217 16289 24281 16353
rect 24297 16289 24361 16353
rect 29637 16289 29701 16353
rect 29717 16289 29781 16353
rect 29797 16289 29861 16353
rect 29877 16289 29941 16353
rect 29957 16289 30021 16353
rect 30037 16289 30101 16353
rect 30117 16289 30181 16353
rect 30197 16289 30261 16353
rect 30277 16289 30341 16353
rect 35643 16297 35707 16361
rect 35723 16297 35787 16361
rect 35803 16297 35867 16361
rect 35883 16297 35947 16361
rect 35963 16297 36027 16361
rect 36043 16297 36107 16361
rect 36123 16297 36187 16361
rect 36203 16297 36267 16361
rect 36283 16297 36347 16361
rect 41639 16285 41703 16349
rect 41719 16285 41783 16349
rect 41799 16285 41863 16349
rect 41879 16285 41943 16349
rect 41959 16285 42023 16349
rect 42039 16285 42103 16349
rect 42119 16285 42183 16349
rect 42199 16285 42263 16349
rect 42279 16285 42343 16349
rect 23635 10958 24339 11102
rect 29629 10950 30333 11094
rect 35599 10938 36303 11082
rect 41627 10962 42331 11106
rect 11663 10530 12367 10674
rect 17633 10550 18337 10694
rect 5640 5224 6344 5368
rect 5652 4842 6356 4986
rect 11648 -337 11712 -273
rect 11728 -337 11792 -273
rect 11808 -337 11872 -273
rect 11888 -337 11952 -273
rect 11968 -337 12032 -273
rect 12048 -337 12112 -273
rect 12128 -337 12192 -273
rect 12208 -337 12272 -273
rect 12288 -337 12352 -273
rect 17636 -325 17700 -261
rect 17716 -325 17780 -261
rect 17796 -325 17860 -261
rect 17876 -325 17940 -261
rect 17956 -325 18020 -261
rect 18036 -325 18100 -261
rect 18116 -325 18180 -261
rect 18196 -325 18260 -261
rect 18276 -325 18340 -261
rect 23745 -766 24449 -622
rect 29807 -786 30511 -642
rect 35651 -766 36355 -622
rect 41653 -774 42357 -630
rect -332 -6003 -268 -5939
rect -252 -6003 -188 -5939
rect -172 -6003 -108 -5939
rect -92 -6003 -28 -5939
rect -12 -6003 52 -5939
rect 68 -6003 132 -5939
rect 148 -6003 212 -5939
rect 228 -6003 292 -5939
rect 5690 -5981 5754 -5917
rect 5770 -5981 5834 -5917
rect 5850 -5981 5914 -5917
rect 5930 -5981 5994 -5917
rect 6010 -5981 6074 -5917
rect 6090 -5981 6154 -5917
rect 6170 -5981 6234 -5917
rect 6250 -5981 6314 -5917
rect 11686 -5991 11750 -5927
rect 11766 -5991 11830 -5927
rect 11846 -5991 11910 -5927
rect 11926 -5991 11990 -5927
rect 12006 -5991 12070 -5927
rect 12086 -5991 12150 -5927
rect 12166 -5991 12230 -5927
rect 12246 -5991 12310 -5927
rect 17686 -5995 17750 -5931
rect 17766 -5995 17830 -5931
rect 17846 -5995 17910 -5931
rect 17926 -5995 17990 -5931
rect 18006 -5995 18070 -5931
rect 18086 -5995 18150 -5931
rect 18166 -5995 18230 -5931
rect 18246 -5995 18310 -5931
rect 23708 -5995 23772 -5931
rect 23788 -5995 23852 -5931
rect 23868 -5995 23932 -5931
rect 23948 -5995 24012 -5931
rect 24028 -5995 24092 -5931
rect 24108 -5995 24172 -5931
rect 24188 -5995 24252 -5931
rect 24268 -5995 24332 -5931
rect 29646 -5987 29710 -5923
rect 29726 -5987 29790 -5923
rect 29806 -5987 29870 -5923
rect 29886 -5987 29950 -5923
rect 29966 -5987 30030 -5923
rect 30046 -5987 30110 -5923
rect 30126 -5987 30190 -5923
rect 30206 -5987 30270 -5923
rect 35686 -5985 35750 -5921
rect 35766 -5985 35830 -5921
rect 35846 -5985 35910 -5921
rect 35926 -5985 35990 -5921
rect 36006 -5985 36070 -5921
rect 36086 -5985 36150 -5921
rect 36166 -5985 36230 -5921
rect 36246 -5985 36310 -5921
rect 41652 -6003 41716 -5939
rect 41732 -6003 41796 -5939
rect 41812 -6003 41876 -5939
rect 41892 -6003 41956 -5939
rect 41972 -6003 42036 -5939
rect 42052 -6003 42116 -5939
rect 42132 -6003 42196 -5939
rect 42212 -6003 42276 -5939
rect -335 -6494 369 -6350
rect 5655 -6464 6359 -6320
rect 11635 -6464 12339 -6320
rect 17639 -6490 18343 -6346
rect 23647 -6464 24351 -6320
rect 29647 -6480 30351 -6336
rect 35631 -6484 36335 -6340
rect 41643 -6468 42347 -6324
rect -922 -17602 -298 -17458
rect 2245 -17604 2949 -17460
rect 8313 -17602 9017 -17458
rect 14263 -17592 14967 -17448
rect 20255 -17588 20959 -17444
rect 26225 -17590 26929 -17446
rect 32245 -17600 32949 -17456
rect 38251 -17594 38955 -17450
rect 44237 -17600 44941 -17456
<< metal4 >>
rect -2130 29562 -1930 29676
rect -3366 29556 -1930 29562
rect -3366 29362 -2460 29556
rect -2130 25094 -1930 29356
rect 10 29332 608 29558
rect 6024 29344 6622 29570
rect 12014 29344 12612 29570
rect 18016 29340 18614 29566
rect 24026 29332 24624 29558
rect 30010 29352 30608 29578
rect 36020 29352 36618 29578
rect 42018 29352 42616 29578
rect 47994 29344 48592 29570
rect -3354 24894 -1930 25094
rect -2130 19428 -1930 24894
rect -3354 19228 -1930 19428
rect -2130 13722 -1930 19228
rect -3366 13522 -1930 13722
rect -2130 8046 -1930 13522
rect -3342 7846 -1930 8046
rect -2130 2340 -1930 7846
rect -3336 2140 -1930 2340
rect -2130 -3294 -1930 2140
rect -3320 -3494 -1930 -3294
rect -2130 -8960 -1930 -3494
rect -3312 -9160 -1930 -8960
rect -2130 -14632 -1930 -9160
rect -3328 -14832 -1930 -14632
rect -2130 -19012 -1930 -14832
rect -702 8198 -498 28418
rect 2184 27982 3018 28020
rect 5292 27998 5496 28018
rect 2184 27838 2283 27982
rect 2907 27838 3018 27982
rect 2184 27798 3018 27838
rect 4970 27937 5828 27998
rect 4970 27873 5056 27937
rect 5120 27873 5136 27937
rect 5200 27873 5216 27937
rect 5280 27873 5296 27937
rect 5360 27873 5376 27937
rect 5440 27873 5456 27937
rect 5520 27873 5536 27937
rect 5600 27873 5616 27937
rect 5680 27873 5696 27937
rect 5760 27873 5828 27937
rect 4970 27798 5828 27873
rect 8204 27978 9038 28012
rect 8204 27834 8289 27978
rect 8913 27834 9038 27978
rect 2 16824 206 27408
rect -396 16756 404 16824
rect -396 16692 -348 16756
rect -284 16692 -268 16756
rect -204 16692 -188 16756
rect -124 16692 -108 16756
rect -44 16692 -28 16756
rect 36 16692 52 16756
rect 116 16692 132 16756
rect 196 16692 212 16756
rect 276 16692 292 16756
rect 356 16692 404 16756
rect -396 16636 404 16692
rect -408 16361 404 16436
rect -408 16297 -351 16361
rect -287 16297 -271 16361
rect -207 16297 -191 16361
rect -127 16297 -111 16361
rect -47 16297 -31 16361
rect 33 16297 49 16361
rect 113 16297 129 16361
rect 193 16297 209 16361
rect 273 16297 289 16361
rect 353 16297 404 16361
rect -408 16224 404 16297
rect -14 11368 202 16224
rect 2530 13570 2730 27798
rect -702 7990 84 8198
rect 5292 8006 5496 27798
rect 8204 27790 9038 27834
rect 14188 27956 15022 28004
rect 14188 27812 14301 27956
rect 14925 27812 15022 27956
rect 5990 16824 6194 27400
rect 5596 16760 6396 16824
rect 5596 16696 5640 16760
rect 5704 16696 5720 16760
rect 5784 16696 5800 16760
rect 5864 16696 5880 16760
rect 5944 16696 5960 16760
rect 6024 16696 6040 16760
rect 6104 16696 6120 16760
rect 6184 16696 6200 16760
rect 6264 16696 6280 16760
rect 6344 16696 6396 16760
rect 5596 16636 6396 16696
rect 5584 16349 6396 16438
rect 5584 16285 5631 16349
rect 5695 16285 5711 16349
rect 5775 16285 5791 16349
rect 5855 16285 5871 16349
rect 5935 16285 5951 16349
rect 6015 16285 6031 16349
rect 6095 16285 6111 16349
rect 6175 16285 6191 16349
rect 6255 16285 6271 16349
rect 6335 16285 6396 16349
rect 5584 16226 6396 16285
rect 5990 11368 6206 16226
rect -702 -17424 -498 7990
rect 4732 7802 5500 8006
rect 8534 7946 8734 27790
rect 14188 27782 15022 27812
rect 20178 27982 21012 28008
rect 20178 27838 20289 27982
rect 20913 27838 21012 27982
rect 20178 27786 21012 27838
rect 26178 27968 27012 28002
rect 26178 27824 26283 27968
rect 26907 27824 27012 27968
rect 11996 16820 12200 27416
rect 11598 16756 12398 16820
rect 11598 16692 11628 16756
rect 11692 16692 11708 16756
rect 11772 16692 11788 16756
rect 11852 16692 11868 16756
rect 11932 16692 11948 16756
rect 12012 16692 12028 16756
rect 12092 16692 12108 16756
rect 12172 16692 12188 16756
rect 12252 16692 12268 16756
rect 12332 16692 12398 16756
rect 11598 16632 12398 16692
rect 11594 16353 12406 16438
rect 11594 16289 11635 16353
rect 11699 16289 11715 16353
rect 11779 16289 11795 16353
rect 11859 16289 11875 16353
rect 11939 16289 11955 16353
rect 12019 16289 12035 16353
rect 12099 16289 12115 16353
rect 12179 16289 12195 16353
rect 12259 16289 12275 16353
rect 12339 16289 12406 16353
rect 11594 16226 12406 16289
rect 11996 11360 12212 16226
rect 11596 10674 12420 10718
rect 11596 10530 11663 10674
rect 12367 10530 12420 10674
rect 11596 10508 12420 10530
rect 4732 7794 5496 7802
rect 4 -5870 210 -1009
rect -410 -5939 398 -5870
rect -410 -6003 -332 -5939
rect -268 -6003 -252 -5939
rect -188 -6003 -172 -5939
rect -108 -6003 -92 -5939
rect -28 -6003 -12 -5939
rect 52 -6003 68 -5939
rect 132 -6003 148 -5939
rect 212 -6003 228 -5939
rect 292 -6003 398 -5939
rect -410 -6064 398 -6003
rect -402 -6350 418 -6312
rect -402 -6494 -335 -6350
rect 369 -6494 418 -6350
rect -402 -6522 418 -6494
rect -10 -17044 210 -6522
rect -1002 -17458 -206 -17424
rect 2534 -17428 2735 2754
rect -1002 -17602 -922 -17458
rect -298 -17602 -206 -17458
rect -1002 -17642 -206 -17602
rect 2198 -17460 3006 -17428
rect 2198 -17604 2245 -17460
rect 2949 -17604 3006 -17460
rect 2198 -17632 3006 -17604
rect -702 -17646 -498 -17642
rect 5292 -18002 5496 7794
rect 5998 5406 6212 6026
rect 12004 5693 12210 10508
rect 14534 7710 14734 27782
rect 17984 16832 18188 27384
rect 17586 16772 18386 16832
rect 17586 16708 17624 16772
rect 17688 16708 17704 16772
rect 17768 16708 17784 16772
rect 17848 16708 17864 16772
rect 17928 16708 17944 16772
rect 18008 16708 18024 16772
rect 18088 16708 18104 16772
rect 18168 16708 18184 16772
rect 18248 16708 18264 16772
rect 18328 16708 18386 16772
rect 17586 16644 18386 16708
rect 17586 16349 18398 16436
rect 17586 16285 17639 16349
rect 17703 16285 17719 16349
rect 17783 16285 17799 16349
rect 17863 16285 17879 16349
rect 17943 16285 17959 16349
rect 18023 16285 18039 16349
rect 18103 16285 18119 16349
rect 18183 16285 18199 16349
rect 18263 16285 18279 16349
rect 18343 16285 18398 16349
rect 17586 16224 18398 16285
rect 18000 11378 18216 16224
rect 17578 10694 18402 10724
rect 17578 10550 17633 10694
rect 18337 10550 18402 10694
rect 17578 10514 18402 10550
rect 17990 5689 18196 10514
rect 20514 7710 20714 27786
rect 26178 27780 27012 27824
rect 32186 27978 33020 28008
rect 32186 27834 32321 27978
rect 32945 27834 33020 27978
rect 32186 27786 33020 27834
rect 38188 27982 39022 28012
rect 38188 27838 38263 27982
rect 38887 27838 39022 27982
rect 38188 27790 39022 27838
rect 44192 27974 45026 28008
rect 44192 27830 44259 27974
rect 44883 27830 45026 27974
rect 23990 16820 24194 27408
rect 23598 16756 24398 16820
rect 23598 16692 23650 16756
rect 23714 16692 23730 16756
rect 23794 16692 23810 16756
rect 23874 16692 23890 16756
rect 23954 16692 23970 16756
rect 24034 16692 24050 16756
rect 24114 16692 24130 16756
rect 24194 16692 24210 16756
rect 24274 16692 24290 16756
rect 24354 16692 24398 16756
rect 23598 16632 24398 16692
rect 23604 16353 24416 16442
rect 23604 16289 23657 16353
rect 23721 16289 23737 16353
rect 23801 16289 23817 16353
rect 23881 16289 23897 16353
rect 23961 16289 23977 16353
rect 24041 16289 24057 16353
rect 24121 16289 24137 16353
rect 24201 16289 24217 16353
rect 24281 16289 24297 16353
rect 24361 16289 24416 16353
rect 23604 16230 24416 16289
rect 24002 11378 24218 16230
rect 23594 11102 24418 11126
rect 23594 10958 23635 11102
rect 24339 10958 24418 11102
rect 23594 10916 24418 10958
rect 23994 5677 24200 10916
rect 26528 7740 26728 27780
rect 29998 16824 30202 27396
rect 29592 16764 30392 16824
rect 29592 16700 29646 16764
rect 29710 16700 29726 16764
rect 29790 16700 29806 16764
rect 29870 16700 29886 16764
rect 29950 16700 29966 16764
rect 30030 16700 30046 16764
rect 30110 16700 30126 16764
rect 30190 16700 30206 16764
rect 30270 16700 30286 16764
rect 30350 16700 30392 16764
rect 29592 16636 30392 16700
rect 29596 16353 30408 16442
rect 29596 16289 29637 16353
rect 29701 16289 29717 16353
rect 29781 16289 29797 16353
rect 29861 16289 29877 16353
rect 29941 16289 29957 16353
rect 30021 16289 30037 16353
rect 30101 16289 30117 16353
rect 30181 16289 30197 16353
rect 30261 16289 30277 16353
rect 30341 16289 30408 16353
rect 29596 16230 30408 16289
rect 29990 11368 30206 16230
rect 29588 11094 30412 11118
rect 29588 10950 29629 11094
rect 30333 10950 30412 11094
rect 29588 10908 30412 10950
rect 30000 5681 30206 10908
rect 32522 7680 32722 27786
rect 35986 16816 36190 27408
rect 35588 16748 36388 16816
rect 35588 16684 35622 16748
rect 35686 16684 35702 16748
rect 35766 16684 35782 16748
rect 35846 16684 35862 16748
rect 35926 16684 35942 16748
rect 36006 16684 36022 16748
rect 36086 16684 36102 16748
rect 36166 16684 36182 16748
rect 36246 16684 36262 16748
rect 36326 16684 36388 16748
rect 35588 16628 36388 16684
rect 35576 16361 36388 16438
rect 35576 16297 35643 16361
rect 35707 16297 35723 16361
rect 35787 16297 35803 16361
rect 35867 16297 35883 16361
rect 35947 16297 35963 16361
rect 36027 16297 36043 16361
rect 36107 16297 36123 16361
rect 36187 16297 36203 16361
rect 36267 16297 36283 16361
rect 36347 16297 36388 16361
rect 35576 16226 36388 16297
rect 35990 11352 36206 16226
rect 35558 11082 36382 11110
rect 35558 10938 35599 11082
rect 36303 10938 36382 11082
rect 35558 10900 36382 10938
rect 35996 5673 36202 10900
rect 38534 7772 38734 27790
rect 44192 27786 45026 27830
rect 41992 16820 42196 27412
rect 41602 16760 42402 16820
rect 41602 16696 41656 16760
rect 41720 16696 41736 16760
rect 41800 16696 41816 16760
rect 41880 16696 41896 16760
rect 41960 16696 41976 16760
rect 42040 16696 42056 16760
rect 42120 16696 42136 16760
rect 42200 16696 42216 16760
rect 42280 16696 42296 16760
rect 42360 16696 42402 16760
rect 41602 16632 42402 16696
rect 41602 16349 42414 16428
rect 41602 16285 41639 16349
rect 41703 16285 41719 16349
rect 41783 16285 41799 16349
rect 41863 16285 41879 16349
rect 41943 16285 41959 16349
rect 42023 16285 42039 16349
rect 42103 16285 42119 16349
rect 42183 16285 42199 16349
rect 42263 16285 42279 16349
rect 42343 16285 42414 16349
rect 41602 16216 42414 16285
rect 41992 11374 42208 16216
rect 41990 11130 42196 11132
rect 41582 11106 42406 11130
rect 41582 10962 41627 11106
rect 42331 10962 42406 11106
rect 41582 10920 42406 10962
rect 41990 5685 42196 10920
rect 44550 7740 44750 27786
rect 49204 25086 49404 29356
rect 48018 24886 49404 25086
rect 49204 19404 49404 24886
rect 47988 19204 49404 19404
rect 49204 13670 49404 19204
rect 47996 13470 49404 13670
rect 49204 8010 49404 13470
rect 48004 7810 49404 8010
rect 5582 5368 6412 5406
rect 5582 5224 5640 5368
rect 6344 5224 6412 5368
rect 5582 5192 6412 5224
rect 5586 4986 6416 5018
rect 5586 4842 5652 4986
rect 6356 4842 6416 4986
rect 5586 4790 6416 4842
rect 5986 4206 6200 4790
rect 5998 -5870 6204 -997
rect 5592 -5917 6400 -5870
rect 5592 -5981 5690 -5917
rect 5754 -5981 5770 -5917
rect 5834 -5981 5850 -5917
rect 5914 -5981 5930 -5917
rect 5994 -5981 6010 -5917
rect 6074 -5981 6090 -5917
rect 6154 -5981 6170 -5917
rect 6234 -5981 6250 -5917
rect 6314 -5981 6400 -5917
rect 5592 -6064 6400 -5981
rect 5604 -6320 6424 -6310
rect 5604 -6464 5655 -6320
rect 6359 -6464 6424 -6320
rect 5604 -6516 6424 -6464
rect 5988 -17020 6208 -6516
rect 8534 -17428 8744 2292
rect 11984 -200 12182 4679
rect 14542 2262 14741 2400
rect 11588 -273 12406 -200
rect 11588 -337 11648 -273
rect 11712 -337 11728 -273
rect 11792 -337 11808 -273
rect 11872 -337 11888 -273
rect 11952 -337 11968 -273
rect 12032 -337 12048 -273
rect 12112 -337 12128 -273
rect 12192 -337 12208 -273
rect 12272 -337 12288 -273
rect 12352 -337 12406 -273
rect 11588 -402 12406 -337
rect 11984 -406 12182 -402
rect 11986 -5870 12192 -993
rect 11592 -5927 12400 -5870
rect 11592 -5991 11686 -5927
rect 11750 -5991 11766 -5927
rect 11830 -5991 11846 -5927
rect 11910 -5991 11926 -5927
rect 11990 -5991 12006 -5927
rect 12070 -5991 12086 -5927
rect 12150 -5991 12166 -5927
rect 12230 -5991 12246 -5927
rect 12310 -5991 12400 -5927
rect 11592 -6064 12400 -5991
rect 11596 -6320 12416 -6302
rect 11596 -6464 11635 -6320
rect 12339 -6464 12416 -6320
rect 11596 -6508 12416 -6464
rect 11994 -17028 12214 -6508
rect 14543 -17428 14740 2262
rect 17996 -196 18194 4679
rect 17600 -261 18418 -196
rect 17600 -325 17636 -261
rect 17700 -325 17716 -261
rect 17780 -325 17796 -261
rect 17860 -325 17876 -261
rect 17940 -325 17956 -261
rect 18020 -325 18036 -261
rect 18100 -325 18116 -261
rect 18180 -325 18196 -261
rect 18260 -325 18276 -261
rect 18340 -325 18418 -261
rect 17600 -398 18418 -325
rect 17986 -5870 18192 -1005
rect 17594 -5931 18402 -5870
rect 17594 -5995 17686 -5931
rect 17750 -5995 17766 -5931
rect 17830 -5995 17846 -5931
rect 17910 -5995 17926 -5931
rect 17990 -5995 18006 -5931
rect 18070 -5995 18086 -5931
rect 18150 -5995 18166 -5931
rect 18230 -5995 18246 -5931
rect 18310 -5995 18402 -5931
rect 17594 -6064 18402 -5995
rect 17588 -6346 18408 -6316
rect 17588 -6490 17639 -6346
rect 18343 -6490 18408 -6346
rect 17588 -6522 18408 -6490
rect 17990 -17024 18210 -6522
rect 20533 -14590 20732 2400
rect 23988 -590 24194 4675
rect 23672 -622 24514 -590
rect 23672 -766 23745 -622
rect 24449 -766 24514 -622
rect 23672 -802 24514 -766
rect 23986 -5870 24192 -997
rect 23586 -5931 24394 -5870
rect 23586 -5995 23708 -5931
rect 23772 -5995 23788 -5931
rect 23852 -5995 23868 -5931
rect 23932 -5995 23948 -5931
rect 24012 -5995 24028 -5931
rect 24092 -5995 24108 -5931
rect 24172 -5995 24188 -5931
rect 24252 -5995 24268 -5931
rect 24332 -5995 24394 -5931
rect 23586 -6064 24394 -5995
rect 23590 -6320 24410 -6302
rect 23590 -6464 23647 -6320
rect 24351 -6464 24410 -6320
rect 23590 -6508 24410 -6464
rect 20532 -14790 20732 -14590
rect 20533 -17424 20732 -14790
rect 23996 -17044 24216 -6508
rect 8240 -17458 9048 -17428
rect 8240 -17602 8313 -17458
rect 9017 -17602 9048 -17458
rect 8240 -17615 9048 -17602
rect 8240 -17632 8534 -17615
rect 8734 -17632 9048 -17615
rect 14200 -17448 15008 -17428
rect 14200 -17592 14263 -17448
rect 14967 -17592 15008 -17448
rect 14200 -17632 15008 -17592
rect 20198 -17444 21006 -17424
rect 26536 -17426 26736 2400
rect 29990 -594 30194 4686
rect 29734 -642 30576 -594
rect 29734 -786 29807 -642
rect 30511 -786 30576 -642
rect 29734 -806 30576 -786
rect 29992 -5874 30198 -993
rect 29544 -5923 30352 -5874
rect 29544 -5987 29646 -5923
rect 29710 -5987 29726 -5923
rect 29790 -5987 29806 -5923
rect 29870 -5987 29886 -5923
rect 29950 -5987 29966 -5923
rect 30030 -5987 30046 -5923
rect 30110 -5987 30126 -5923
rect 30190 -5987 30206 -5923
rect 30270 -5987 30352 -5923
rect 29544 -6068 30352 -5987
rect 29594 -6336 30414 -6310
rect 29594 -6480 29647 -6336
rect 30351 -6480 30414 -6336
rect 29594 -6516 30414 -6480
rect 29996 -17036 30216 -6516
rect 20198 -17588 20255 -17444
rect 20959 -17588 21006 -17444
rect 20198 -17628 21006 -17588
rect 26192 -17446 27000 -17426
rect 32532 -17430 32732 2400
rect 35992 -590 36196 4678
rect 35610 -622 36420 -590
rect 35610 -766 35651 -622
rect 36355 -766 36420 -622
rect 35610 -798 36420 -766
rect 35996 -5870 36202 -997
rect 35578 -5921 36386 -5870
rect 35578 -5985 35686 -5921
rect 35750 -5985 35766 -5921
rect 35830 -5985 35846 -5921
rect 35910 -5985 35926 -5921
rect 35990 -5985 36006 -5921
rect 36070 -5985 36086 -5921
rect 36150 -5985 36166 -5921
rect 36230 -5985 36246 -5921
rect 36310 -5985 36386 -5921
rect 35578 -6064 36386 -5985
rect 35584 -6340 36404 -6302
rect 35584 -6484 35631 -6340
rect 36335 -6484 36404 -6340
rect 35584 -6508 36404 -6484
rect 35996 -17028 36216 -6508
rect 38536 -17430 38736 2400
rect 41990 -590 42194 4686
rect 41596 -630 42406 -590
rect 41596 -774 41653 -630
rect 42357 -774 42406 -630
rect 41596 -798 42406 -774
rect 41982 -5874 42188 -1013
rect 41576 -5939 42384 -5874
rect 41576 -6003 41652 -5939
rect 41716 -6003 41732 -5939
rect 41796 -6003 41812 -5939
rect 41876 -6003 41892 -5939
rect 41956 -6003 41972 -5939
rect 42036 -6003 42052 -5939
rect 42116 -6003 42132 -5939
rect 42196 -6003 42212 -5939
rect 42276 -6003 42384 -5939
rect 41576 -6068 42384 -6003
rect 41588 -6324 42408 -6302
rect 41588 -6468 41643 -6324
rect 42347 -6468 42408 -6324
rect 41588 -6508 42408 -6468
rect 41994 -17020 42214 -6508
rect 44510 -17426 44710 2400
rect 49204 2322 49404 7810
rect 47988 2122 49404 2322
rect 49204 -3284 49404 2122
rect 48026 -3484 49404 -3284
rect 49204 -8928 49404 -3484
rect 48004 -9128 49404 -8928
rect 49204 -14732 49404 -9128
rect 48042 -14932 49404 -14732
rect 26192 -17590 26225 -17446
rect 26929 -17590 27000 -17446
rect 20533 -17631 20732 -17628
rect 26192 -17630 27000 -17590
rect 32194 -17456 33002 -17430
rect 32194 -17600 32245 -17456
rect 32949 -17600 33002 -17456
rect 26536 -17632 26736 -17630
rect 14543 -17642 14740 -17632
rect 32194 -17634 33002 -17600
rect 38196 -17450 39004 -17430
rect 38196 -17594 38251 -17450
rect 38955 -17594 39004 -17450
rect 38196 -17634 39004 -17594
rect 44196 -17456 45004 -17426
rect 44196 -17600 44237 -17456
rect 44941 -17600 45004 -17456
rect 44196 -17630 45004 -17600
rect 32532 -17636 32732 -17634
rect 38536 -17642 38736 -17634
rect -3346 -19212 -1022 -19012
rect -26 -19214 572 -18988
rect 5992 -19218 6590 -18992
rect 11998 -19210 12596 -18984
rect 17998 -19210 18596 -18984
rect 24008 -19198 24606 -18972
rect 30018 -19198 30616 -18972
rect 36016 -19210 36614 -18984
rect 42010 -19194 42608 -18968
rect 49204 -19044 49404 -14932
rect 48014 -19244 49404 -19044
rect 48018 -19280 49404 -19244
use core1r  core1r_0
timestamp 1699926577
transform 1 0 0 0 1 -11356
box 0 0 46972 4680
use core1r  core1r_1
timestamp 1699926577
transform 1 0 0 0 1 -5680
box 0 0 46972 4680
use core1r  core1r_2
timestamp 1699926577
transform 1 0 0 0 1 22720
box 0 0 46972 4680
use core1r  core1r_3
timestamp 1699926577
transform 1 0 0 0 1 -17036
box 0 0 46972 4680
use core1r  core1r_4
timestamp 1699926577
transform 1 0 0 0 1 11360
box 0 0 46972 4680
use core1r  core1r_5
timestamp 1699926577
transform 1 0 0 0 1 17040
box 0 0 46972 4680
use core2r  core2r_0
timestamp 1699926577
transform 1 0 0 0 1 5680
box 0 -5680 46972 4680
use d1rleftright  d1rleftright_0
timestamp 1699926577
transform 1 0 47976 0 1 -17032
box 0 0 2372 44440
use d1rleftright  d1rleftright_1
timestamp 1699926577
transform 1 0 -3374 0 1 -17036
box 0 0 2372 44440
use d1rtopbottom  d1rtopbottom_0
timestamp 1699926577
transform 1 0 0 0 1 -20114
box 0 0 46972 2080
use d1rtopbottom  d1rtopbottom_1
timestamp 1699926577
transform 1 0 0 0 1 28400
box 0 0 46972 2080
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_0
timestamp 1699926577
transform -1 0 49158 0 1 29440
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_1
timestamp 1699926577
transform -1 0 49158 0 1 -19074
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_2
timestamp 1699926577
transform -1 0 -2186 0 1 -19078
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_3
timestamp 1699926577
transform -1 0 -2188 0 1 29444
box -1186 -1040 1186 1040
<< labels >>
flabel metal3 s -3422 4806 -2566 5002 0 FreeSans 6326 0 0 0 D0
port 1 nsew
flabel metal3 s -3408 5214 -2552 5410 0 FreeSans 6326 0 0 0 D5
port 2 nsew
flabel metal3 s -3406 -400 -2580 -200 0 FreeSans 6326 0 0 0 D1
port 3 nsew
flabel metal3 s -3414 -796 -2588 -596 0 FreeSans 6326 0 0 0 D2
port 4 nsew
flabel metal3 s -3208 -6050 -2386 -5878 0 FreeSans 6326 0 0 0 D3
port 5 nsew
flabel metal3 s -3192 -6506 -2370 -6334 0 FreeSans 6326 0 0 0 D4
port 6 nsew
flabel metal3 s -3214 10524 -2390 10734 0 FreeSans 6326 0 0 0 D6
port 7 nsew
flabel metal3 s -3194 10920 -2370 11130 0 FreeSans 6326 0 0 0 D7
port 8 nsew
flabel metal3 s -3192 16230 -2380 16442 0 FreeSans 6326 0 0 0 D8
port 9 nsew
flabel metal3 s -3198 16624 -2386 16836 0 FreeSans 6326 0 0 0 D9
port 10 nsew
flabel metal4 s -702 7990 -314 8190 0 FreeSans 6326 0 0 0 VP1
port 11 nsew
flabel metal4 s 5216 7802 5500 8006 0 FreeSans 6326 0 0 0 VP2
port 12 nsew
flabel metal3 s 5142 -19198 5782 -18970 0 FreeSans 6326 0 0 0 VSS
port 13 nsew
<< end >>
