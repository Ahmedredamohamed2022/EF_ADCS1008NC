VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO EF_ADCS1008NC
  CLASS BLOCK ;
  FOREIGN EF_ADCS1008NC ;
  ORIGIN 0.000 0.000 ;
  SIZE 344.540 BY 524.120 ;
  PIN HOLD
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.360000 ;
    PORT
      LAYER met3 ;
        RECT 0.680 439.985 3.880 440.995 ;
    END
    PORT
      LAYER met1 ;
        RECT 6.550 439.970 7.550 440.970 ;
    END
  END HOLD
  PIN EN
    ANTENNAGATEAREA 1.752000 ;
    ANTENNADIFFAREA 1.080000 ;
    PORT
      LAYER met3 ;
        RECT 0.680 418.755 3.480 419.685 ;
    END
  END EN
  PIN RST
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER met3 ;
        RECT 0.680 383.285 3.180 384.295 ;
    END
  END RST
  PIN DATA[9]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.680 325.735 3.450 326.615 ;
    END
  END DATA[9]
  PIN DATA[8]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.680 292.105 3.920 292.985 ;
    END
  END DATA[8]
  PIN DATA[7]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.680 258.525 3.920 259.405 ;
    END
  END DATA[7]
  PIN DATA[6]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.680 225.055 3.920 225.935 ;
    END
  END DATA[6]
  PIN DATA[5]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.680 191.205 3.920 192.085 ;
    END
  END DATA[5]
  PIN DATA[0]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.680 156.275 3.920 157.155 ;
    END
  END DATA[0]
  PIN DATA[1]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.680 122.745 3.920 123.625 ;
    END
  END DATA[1]
  PIN DATA[2]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.680 89.145 3.920 90.025 ;
    END
  END DATA[2]
  PIN DATA[3]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.680 55.635 3.920 56.515 ;
    END
  END DATA[3]
  PIN DATA[4]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.680 21.745 3.920 22.625 ;
    END
  END DATA[4]
  PIN DVSS
    ANTENNAGATEAREA 74.759102 ;
    ANTENNADIFFAREA 1023.766663 ;
    PORT
      LAYER met3 ;
        RECT 0.680 11.375 5.120 13.375 ;
    END
  END DVSS
  PIN DVDD
    ANTENNAGATEAREA 47.261497 ;
    ANTENNADIFFAREA 93.596451 ;
    PORT
      LAYER met3 ;
        RECT 0.680 14.055 5.120 16.055 ;
    END
  END DVDD
  PIN VDD
    ANTENNAGATEAREA 100.000000 ;
    ANTENNADIFFAREA 2509.495605 ;
    PORT
      LAYER met3 ;
        RECT 0.680 8.915 5.300 10.875 ;
    END
  END VDD
  PIN VH
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met3 ;
        RECT 0.680 186.645 3.970 187.525 ;
    END
  END VH
  PIN VL
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met3 ;
        RECT 0.680 184.315 3.970 185.195 ;
    END
  END VL
  PIN VSS
    ANTENNAGATEAREA 130.500000 ;
    ANTENNADIFFAREA 621.362671 ;
    PORT
      LAYER met3 ;
        RECT 0.680 6.120 6.800 8.050 ;
    END
  END VSS
  PIN CMP
    ANTENNADIFFAREA 0.492900 ;
    PORT
      LAYER met2 ;
        RECT 182.680 522.150 183.670 524.110 ;
    END
  END CMP
  PIN VIN[7]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 22.800 522.270 23.270 524.120 ;
    END
  END VIN[7]
  PIN VIN[6]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 39.820 522.270 40.290 524.120 ;
    END
  END VIN[6]
  PIN VIN[5]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 56.810 522.270 57.280 524.120 ;
    END
  END VIN[5]
  PIN VIN[4]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 73.320 522.270 73.790 524.120 ;
    END
  END VIN[4]
  PIN VIN[3]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 89.880 522.270 90.350 524.120 ;
    END
  END VIN[3]
  PIN VIN[2]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 106.740 522.270 107.210 524.120 ;
    END
  END VIN[2]
  PIN VIN[1]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 123.250 522.270 123.720 524.120 ;
    END
  END VIN[1]
  PIN VIN[0]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 140.480 522.270 140.950 524.120 ;
    END
  END VIN[0]
  PIN B[0]
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 176.630 522.120 176.980 524.120 ;
    END
  END B[0]
  PIN B[1]
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 177.360 522.120 177.710 524.120 ;
    END
  END B[1]
  PIN B[2]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 178.090 522.120 178.440 524.120 ;
    END
  END B[2]
  OBS
      LAYER li1 ;
        RECT 7.455 20.205 248.590 513.925 ;
      LAYER met1 ;
        RECT 0.735 441.250 249.285 514.130 ;
        RECT 0.735 439.690 6.270 441.250 ;
        RECT 7.830 439.690 249.285 441.250 ;
        RECT 0.735 17.890 249.285 439.690 ;
      LAYER met2 ;
        RECT 0.690 521.990 22.520 524.120 ;
        RECT 23.550 521.990 39.540 524.120 ;
        RECT 40.570 521.990 56.530 524.120 ;
        RECT 57.560 521.990 73.040 524.120 ;
        RECT 74.070 521.990 89.600 524.120 ;
        RECT 90.630 521.990 106.460 524.120 ;
        RECT 107.490 521.990 122.970 524.120 ;
        RECT 124.000 521.990 140.200 524.120 ;
        RECT 141.230 521.990 176.350 524.120 ;
        RECT 0.690 521.840 176.350 521.990 ;
        RECT 178.720 521.870 182.400 524.120 ;
        RECT 183.950 521.870 246.970 524.120 ;
        RECT 178.720 521.840 246.970 521.870 ;
        RECT 0.690 17.890 246.970 521.840 ;
      LAYER met3 ;
        RECT 0.680 441.395 344.540 523.970 ;
        RECT 4.280 439.585 344.540 441.395 ;
        RECT 0.680 420.085 344.540 439.585 ;
        RECT 3.880 418.355 344.540 420.085 ;
        RECT 0.680 384.695 344.540 418.355 ;
        RECT 3.580 382.885 344.540 384.695 ;
        RECT 0.680 327.015 344.540 382.885 ;
        RECT 3.850 325.335 344.540 327.015 ;
        RECT 0.680 293.385 344.540 325.335 ;
        RECT 4.320 291.705 344.540 293.385 ;
        RECT 0.680 259.805 344.540 291.705 ;
        RECT 4.320 258.125 344.540 259.805 ;
        RECT 0.680 226.335 344.540 258.125 ;
        RECT 4.320 224.655 344.540 226.335 ;
        RECT 0.680 192.485 344.540 224.655 ;
        RECT 4.320 190.805 344.540 192.485 ;
        RECT 0.680 187.925 344.540 190.805 ;
        RECT 4.370 186.245 344.540 187.925 ;
        RECT 0.680 185.595 344.540 186.245 ;
        RECT 4.370 183.915 344.540 185.595 ;
        RECT 0.680 157.555 344.540 183.915 ;
        RECT 4.320 155.875 344.540 157.555 ;
        RECT 0.680 124.025 344.540 155.875 ;
        RECT 4.320 122.345 344.540 124.025 ;
        RECT 0.680 90.425 344.540 122.345 ;
        RECT 4.320 88.745 344.540 90.425 ;
        RECT 0.680 56.915 344.540 88.745 ;
        RECT 4.320 55.235 344.540 56.915 ;
        RECT 0.680 23.025 344.540 55.235 ;
        RECT 4.320 21.345 344.540 23.025 ;
        RECT 0.680 16.455 344.540 21.345 ;
        RECT 5.520 11.275 344.540 16.455 ;
        RECT 5.700 8.515 344.540 11.275 ;
        RECT 0.680 8.450 344.540 8.515 ;
        RECT 7.200 6.120 344.540 8.450 ;
      LAYER met4 ;
        RECT 4.560 6.130 344.370 521.730 ;
      LAYER met5 ;
        RECT 17.165 390.585 171.645 512.900 ;
  END
END EF_ADCS1008NC
END LIBRARY

