magic
tech sky130A
magscale 1 2
timestamp 1699926577
<< pwell >>
rect -188 -188 188 188
<< psubdiff >>
rect -162 128 -51 162
rect -17 128 17 162
rect 51 128 162 162
rect -162 51 -128 128
rect -162 -17 -128 17
rect -162 -128 -128 -51
rect 128 51 162 128
rect 128 -17 162 17
rect 128 -128 162 -51
rect -162 -162 -51 -128
rect -17 -162 17 -128
rect 51 -162 162 -128
<< psubdiffcont >>
rect -51 128 -17 162
rect 17 128 51 162
rect -162 17 -128 51
rect -162 -51 -128 -17
rect 128 17 162 51
rect 128 -51 162 -17
rect -51 -162 -17 -128
rect 17 -162 51 -128
<< ndiode >>
rect -60 17 60 60
rect -60 -17 -17 17
rect 17 -17 60 17
rect -60 -60 60 -17
<< ndiodec >>
rect -17 -17 17 17
<< locali >>
rect -162 128 -51 162
rect -17 128 17 162
rect 51 128 162 162
rect -162 51 -128 128
rect 128 51 162 128
rect -162 -17 -128 17
rect -64 17 64 48
rect -64 -17 -17 17
rect 17 -17 64 17
rect -64 -48 64 -17
rect 128 -17 162 17
rect -162 -128 -128 -51
rect 128 -128 162 -51
rect -162 -162 -51 -128
rect -17 -162 17 -128
rect 51 -162 162 -128
<< viali >>
rect -17 -17 17 17
<< metal1 >>
rect -60 17 60 54
rect -60 -17 -17 17
rect 17 -17 60 17
rect -60 -54 60 -17
<< properties >>
string FIXED_BBOX -144 -144 144 144
<< end >>
