magic
tech sky130A
magscale 1 2
timestamp 1699926577
<< metal1 >>
rect 21620 68923 21824 68936
rect 21617 68888 21824 68923
rect 21617 68388 21664 68888
rect 21780 68388 21824 68888
rect 21617 68344 21824 68388
rect 10320 60008 10452 60010
rect 8076 59993 10452 60008
rect 8076 59941 10355 59993
rect 10407 59941 10452 59993
rect 8076 59929 10452 59941
rect 8076 59877 10355 59929
rect 10407 59877 10452 59929
rect 8076 59865 10452 59877
rect 8076 59813 10355 59865
rect 10407 59813 10452 59865
rect 8076 59790 10452 59813
rect 8076 59786 10446 59790
rect 17156 57056 17362 57256
rect 17156 56951 17358 57056
rect 21617 56951 21819 68344
rect 26976 66578 27604 68210
rect 26976 66142 27041 66578
rect 27541 66142 27604 66578
rect 26976 59544 27604 66142
rect 33784 67395 34206 68225
rect 33784 66895 33836 67395
rect 34144 66895 34206 67395
rect 33784 62990 34206 66895
rect 35986 68112 36420 68190
rect 35986 67676 36046 68112
rect 36354 67676 36420 68112
rect 35986 62700 36420 67676
rect 35986 62392 36043 62700
rect 36351 62392 36420 62700
rect 35986 62354 36420 62392
rect 26976 59044 27036 59544
rect 27536 59044 27604 59544
rect 26976 58990 27604 59044
rect 1362 56460 1480 56776
rect 17156 56749 21819 56951
rect 28358 55812 28550 58174
rect 28002 55774 28856 55812
rect 28002 55658 28034 55774
rect 28790 55658 28856 55774
rect 28002 55604 28856 55658
rect 31654 55426 31846 58072
rect 43194 57198 43376 57612
rect 43188 57190 43990 57198
rect 41915 57162 43990 57190
rect 41915 57046 43256 57162
rect 43948 57046 43990 57162
rect 41915 57020 43990 57046
rect 43188 57008 43990 57020
rect 42396 55426 43234 55434
rect 10758 55400 47567 55426
rect 10758 55220 13014 55400
rect 13642 55376 47567 55400
rect 13642 55375 42453 55376
rect 13642 55259 31220 55375
rect 32104 55260 42453 55375
rect 43209 55260 47567 55376
rect 32104 55259 47567 55260
rect 13642 55220 47567 55259
rect 12984 55216 13684 55220
rect 12988 55202 13682 55216
rect 31202 55194 32136 55220
rect 42396 55212 43234 55220
rect 10118 53244 10236 53256
rect 8042 53238 10440 53244
rect 8042 53186 10152 53238
rect 10204 53186 10440 53238
rect 8042 53174 10440 53186
rect 8042 53122 10152 53174
rect 10204 53122 10440 53174
rect 8042 53110 10440 53122
rect 8042 53058 10152 53110
rect 10204 53058 10440 53110
rect 8042 53026 10440 53058
rect 1342 49738 1460 50054
rect 7994 46503 10436 46518
rect 7994 46451 9964 46503
rect 10016 46451 10436 46503
rect 7994 46439 10436 46451
rect 7994 46387 9964 46439
rect 10016 46387 10436 46439
rect 7994 46375 10436 46387
rect 7994 46323 9964 46375
rect 10016 46323 10436 46375
rect 7994 46310 10436 46323
rect 9912 46304 10050 46310
rect 1342 43020 1460 43336
rect 8156 39790 10446 39810
rect 8156 39738 9764 39790
rect 9816 39738 10446 39790
rect 8156 39726 10446 39738
rect 8156 39674 9764 39726
rect 9816 39674 10446 39726
rect 8156 39662 10446 39674
rect 8156 39610 9764 39662
rect 9816 39610 10446 39662
rect 8156 39600 10446 39610
rect 8152 39592 10446 39600
rect 9728 39588 9854 39592
rect 1334 36334 1452 36650
rect 8060 32990 10436 33010
rect 8060 32938 9541 32990
rect 9593 32938 10436 32990
rect 8060 32926 10436 32938
rect 8060 32874 9541 32926
rect 9593 32874 10436 32926
rect 8060 32862 10436 32874
rect 8060 32810 9541 32862
rect 9593 32810 10436 32862
rect 8060 32790 10436 32810
rect 1348 29550 1466 29866
rect 8060 26062 10436 26072
rect 8060 26010 8522 26062
rect 8574 26010 10436 26062
rect 8060 25998 10436 26010
rect 8060 25946 8522 25998
rect 8574 25946 10436 25998
rect 8060 25934 10436 25946
rect 8060 25882 8522 25934
rect 8574 25882 10436 25934
rect 8060 25868 10436 25882
rect 8488 25864 8604 25868
rect 1356 22592 1474 22908
rect 8690 19400 8812 19406
rect 8002 19370 10434 19400
rect 8002 19318 8726 19370
rect 8778 19318 10434 19370
rect 8002 19306 10434 19318
rect 8002 19254 8726 19306
rect 8778 19254 10434 19306
rect 8002 19204 10434 19254
rect 1350 15862 1468 16178
rect 8058 12557 10438 12600
rect 8058 12505 8920 12557
rect 8972 12505 10438 12557
rect 8058 12493 10438 12505
rect 8058 12441 8920 12493
rect 8972 12441 10438 12493
rect 8058 12396 10438 12441
rect 8890 12394 9008 12396
rect 1342 9144 1460 9460
rect 7990 5960 10436 6002
rect 7990 5908 9122 5960
rect 9174 5908 10436 5960
rect 7990 5896 10436 5908
rect 7990 5844 9122 5896
rect 9174 5844 10436 5896
rect 7990 5798 10436 5844
rect 1330 2452 1448 2768
rect 9298 -792 9416 -786
rect 8064 -811 10432 -792
rect 8064 -863 9333 -811
rect 9385 -863 10432 -811
rect 8064 -875 10432 -863
rect 8064 -927 9333 -875
rect 9385 -927 10432 -875
rect 8064 -939 10432 -927
rect 8064 -991 9333 -939
rect 9385 -991 10432 -939
rect 8064 -1006 10432 -991
rect 9298 -1012 9416 -1006
rect 1328 -4080 1464 -3984
rect 1328 -4338 1464 -4306
rect 1750 -4414 2216 -4374
rect 1750 -4658 1811 -4414
rect 2183 -4658 2216 -4414
rect 1750 -4738 2216 -4658
<< via1 >>
rect 21664 68388 21780 68888
rect 10355 59941 10407 59993
rect 10355 59877 10407 59929
rect 10355 59813 10407 59865
rect 27041 66142 27541 66578
rect 33836 66895 34144 67395
rect 36046 67676 36354 68112
rect 36043 62392 36351 62700
rect 27036 59044 27536 59544
rect 28034 55658 28790 55774
rect 43256 57046 43948 57162
rect 13014 55220 13642 55400
rect 31220 55259 32104 55375
rect 42453 55260 43209 55376
rect 10152 53186 10204 53238
rect 10152 53122 10204 53174
rect 10152 53058 10204 53110
rect 9964 46451 10016 46503
rect 9964 46387 10016 46439
rect 9964 46323 10016 46375
rect 9764 39738 9816 39790
rect 9764 39674 9816 39726
rect 9764 39610 9816 39662
rect 9541 32938 9593 32990
rect 9541 32874 9593 32926
rect 9541 32810 9593 32862
rect 8522 26010 8574 26062
rect 8522 25946 8574 25998
rect 8522 25882 8574 25934
rect 8726 19318 8778 19370
rect 8726 19254 8778 19306
rect 8920 12505 8972 12557
rect 8920 12441 8972 12493
rect 9122 5908 9174 5960
rect 9122 5844 9174 5896
rect 9333 -863 9385 -811
rect 9333 -927 9385 -875
rect 9333 -991 9385 -939
rect 1811 -4658 2183 -4414
<< metal2 >>
rect 17206 68986 17426 68998
rect 17200 68976 17432 68986
rect 17200 68318 17448 68976
rect 21620 68888 21824 68936
rect 21620 68388 21664 68888
rect 21780 68388 21824 68888
rect 21620 68344 21824 68388
rect 17206 68308 17448 68318
rect 17228 67794 17448 68308
rect 30190 68212 30412 68814
rect 17200 66764 17448 67794
rect 17228 64992 17448 66764
rect 26994 66578 27586 66616
rect 26994 66142 27041 66578
rect 27541 66142 27586 66578
rect 26994 66042 27586 66142
rect 17212 64632 17448 64992
rect 17228 64018 17448 64632
rect 30196 63508 30412 68212
rect 35992 68122 36410 68178
rect 35992 68112 36052 68122
rect 36348 68112 36410 68122
rect 35992 67676 36046 68112
rect 36354 67676 36410 68112
rect 35992 67666 36052 67676
rect 36348 67666 36410 67676
rect 35992 67610 36410 67666
rect 33776 67395 34206 67436
rect 33776 66895 33836 67395
rect 34144 66895 34206 67395
rect 33776 66826 34206 66895
rect 29724 63435 31084 63508
rect 29724 63299 29796 63435
rect 31052 63299 31084 63435
rect 29724 63252 31084 63299
rect 35992 62700 36416 62776
rect 35992 62392 36043 62700
rect 36351 62392 36416 62700
rect 35992 62330 36416 62392
rect 10320 59993 10452 60010
rect 10320 59971 10355 59993
rect 10407 59971 10452 59993
rect 10320 59915 10353 59971
rect 10409 59915 10452 59971
rect 10320 59891 10355 59915
rect 10407 59891 10452 59915
rect 10320 59835 10353 59891
rect 10409 59835 10452 59891
rect 10320 59813 10355 59835
rect 10407 59813 10452 59835
rect 10320 59790 10452 59813
rect 26976 59544 27622 59608
rect 26976 59044 27036 59544
rect 27536 59044 27622 59544
rect 26976 58990 27622 59044
rect 41874 57585 42618 57602
rect 15380 57365 16564 57404
rect 15380 57229 15411 57365
rect 16507 57229 16564 57365
rect 15380 57188 16564 57229
rect -400 56949 1908 57003
rect -400 56893 -377 56949
rect -321 56893 -297 56949
rect -241 56893 -217 56949
rect -161 56893 -137 56949
rect -81 56893 -57 56949
rect -1 56893 23 56949
rect 79 56893 103 56949
rect 159 56893 1908 56949
rect -400 56831 1908 56893
rect 16816 56598 17018 57454
rect 41874 57449 41898 57585
rect 42594 57449 42618 57585
rect 41874 57432 42618 57449
rect 17616 57316 18796 57320
rect 17616 57180 17618 57316
rect 18794 57180 18796 57316
rect 17616 57176 18796 57180
rect 42846 56654 43012 57735
rect 43578 57198 43982 57626
rect 43188 57171 43990 57198
rect 43188 57035 43234 57171
rect 43930 57162 43990 57171
rect 43948 57046 43990 57162
rect 43930 57035 43990 57046
rect 43188 57008 43990 57035
rect 43578 57004 43982 57008
rect 16796 56388 17020 56598
rect 42820 56444 43044 56654
rect 16816 55816 17018 56388
rect 16542 55775 17336 55816
rect 16542 55639 16584 55775
rect 17280 55639 17336 55775
rect 16542 55596 17336 55639
rect 28002 55784 28856 55812
rect 28002 55648 28024 55784
rect 28800 55648 28856 55784
rect 28002 55604 28856 55648
rect 16816 55595 17018 55596
rect 42846 55434 43012 56444
rect 12988 55408 13682 55420
rect 12984 55400 13684 55408
rect 42396 55406 43234 55434
rect 12984 55220 13014 55400
rect 13642 55220 13684 55400
rect 12984 55216 13684 55220
rect 31202 55375 32136 55406
rect 31202 55259 31220 55375
rect 32104 55259 32136 55375
rect 12988 55202 13682 55216
rect 31202 55194 32136 55259
rect 42394 55376 43242 55406
rect 42394 55260 42453 55376
rect 43209 55260 43242 55376
rect 42394 55190 43242 55260
rect 42846 55189 43012 55190
rect 10118 53238 10236 53256
rect 10118 53216 10152 53238
rect 10204 53216 10236 53238
rect 10118 53160 10150 53216
rect 10206 53160 10236 53216
rect 10118 53136 10152 53160
rect 10204 53136 10236 53160
rect 10118 53080 10150 53136
rect 10206 53080 10236 53136
rect 10118 53058 10152 53080
rect 10204 53058 10236 53080
rect 10118 53038 10236 53058
rect -402 50264 1882 50275
rect -402 50128 -364 50264
rect 172 50128 1882 50264
rect -402 50103 1882 50128
rect 9912 46503 10050 46512
rect 9912 46481 9964 46503
rect 10016 46481 10050 46503
rect 9912 46425 9962 46481
rect 10018 46425 10050 46481
rect 9912 46401 9964 46425
rect 10016 46401 10050 46425
rect 9912 46345 9962 46401
rect 10018 46345 10050 46401
rect 9912 46323 9964 46345
rect 10016 46323 10050 46345
rect 9912 46304 10050 46323
rect -400 43503 1880 43561
rect -400 43447 -378 43503
rect -322 43447 -298 43503
rect -242 43447 -218 43503
rect -162 43447 -138 43503
rect -82 43447 -58 43503
rect -2 43447 22 43503
rect 78 43447 102 43503
rect 158 43447 1880 43503
rect -400 43389 1880 43447
rect 9728 39790 9854 39804
rect 9728 39768 9764 39790
rect 9816 39768 9854 39790
rect 9728 39712 9762 39768
rect 9818 39712 9854 39768
rect 9728 39688 9764 39712
rect 9816 39688 9854 39712
rect 9728 39632 9762 39688
rect 9818 39632 9854 39688
rect 9728 39610 9764 39632
rect 9816 39610 9854 39632
rect 9728 39588 9854 39610
rect -400 36860 1882 36871
rect -400 36724 -377 36860
rect 159 36724 1882 36860
rect -400 36699 1882 36724
rect 9502 32990 9632 33008
rect 9502 32968 9541 32990
rect 9593 32968 9632 32990
rect 9502 32912 9539 32968
rect 9595 32912 9632 32968
rect 9502 32888 9541 32912
rect 9593 32888 9632 32912
rect 9502 32832 9539 32888
rect 9595 32832 9632 32888
rect 9502 32810 9541 32832
rect 9593 32810 9632 32832
rect 9502 32790 9632 32810
rect -406 30077 1804 30089
rect -406 29941 -379 30077
rect 157 29941 1804 30077
rect -406 29917 1804 29941
rect 8488 26062 8604 26070
rect 8488 26040 8522 26062
rect 8574 26040 8604 26062
rect 8488 25984 8520 26040
rect 8576 25984 8604 26040
rect 8488 25960 8522 25984
rect 8574 25960 8604 25984
rect 8488 25904 8520 25960
rect 8576 25904 8604 25960
rect 8488 25882 8522 25904
rect 8574 25882 8604 25904
rect 8488 25864 8604 25882
rect -402 23071 1908 23119
rect -402 23015 -364 23071
rect -308 23015 -284 23071
rect -228 23015 -204 23071
rect -148 23015 -124 23071
rect -68 23015 -44 23071
rect 12 23015 36 23071
rect 92 23015 116 23071
rect 172 23015 1908 23071
rect -402 22947 1908 23015
rect 8690 19380 8812 19406
rect 8690 19324 8724 19380
rect 8780 19324 8812 19380
rect 8690 19318 8726 19324
rect 8778 19318 8812 19324
rect 8690 19306 8812 19318
rect 8690 19300 8726 19306
rect 8778 19300 8812 19306
rect 8690 19244 8724 19300
rect 8780 19244 8812 19300
rect 8690 19210 8812 19244
rect -400 16337 1866 16391
rect -400 16281 -376 16337
rect -320 16281 -296 16337
rect -240 16281 -216 16337
rect -160 16281 -136 16337
rect -80 16281 -56 16337
rect 0 16281 24 16337
rect 80 16281 104 16337
rect 160 16281 1866 16337
rect -400 16219 1866 16281
rect 8890 12567 9008 12598
rect 8890 12511 8918 12567
rect 8974 12511 9008 12567
rect 8890 12505 8920 12511
rect 8972 12505 9008 12511
rect 8890 12493 9008 12505
rect 8890 12487 8920 12493
rect 8972 12487 9008 12493
rect 8890 12431 8918 12487
rect 8974 12431 9008 12487
rect 8890 12394 9008 12431
rect -402 9634 1870 9677
rect -402 9578 -374 9634
rect -318 9578 -294 9634
rect -238 9578 -214 9634
rect -158 9578 -134 9634
rect -78 9578 -54 9634
rect 2 9578 26 9634
rect 82 9578 106 9634
rect 162 9578 1870 9634
rect -402 9505 1870 9578
rect 9086 5970 9200 6002
rect 9086 5914 9120 5970
rect 9176 5914 9200 5970
rect 9086 5908 9122 5914
rect 9174 5908 9200 5914
rect 9086 5896 9200 5908
rect 9086 5890 9122 5896
rect 9174 5890 9200 5896
rect 9086 5834 9120 5890
rect 9176 5834 9200 5890
rect 9086 5798 9200 5834
rect -402 2980 1794 2987
rect -402 2844 -380 2980
rect 156 2844 1794 2980
rect -402 2815 1794 2844
rect 9298 -811 9416 -786
rect 9298 -833 9333 -811
rect 9385 -833 9416 -811
rect 9298 -889 9331 -833
rect 9387 -889 9416 -833
rect 9298 -913 9333 -889
rect 9385 -913 9416 -889
rect 9298 -969 9331 -913
rect 9387 -969 9416 -913
rect 9298 -991 9333 -969
rect 9385 -991 9416 -969
rect 9298 -1012 9416 -991
rect -400 -3814 1896 -3795
rect -400 -3950 -377 -3814
rect 159 -3950 1896 -3814
rect -400 -3967 1896 -3950
rect 1750 -4414 2216 -4374
rect 1750 -4428 1811 -4414
rect 2183 -4428 2216 -4414
rect 1750 -4644 1809 -4428
rect 2185 -4644 2216 -4428
rect 1750 -4658 1811 -4644
rect 2183 -4658 2216 -4644
rect 1750 -4738 2216 -4658
<< via2 >>
rect 27063 66172 27519 66548
rect 36052 68112 36348 68122
rect 36052 67676 36348 68112
rect 36052 67666 36348 67676
rect 33842 66917 34138 67373
rect 29796 63299 31052 63435
rect 36049 62398 36345 62694
rect 10353 59941 10355 59971
rect 10355 59941 10407 59971
rect 10407 59941 10409 59971
rect 10353 59929 10409 59941
rect 10353 59915 10355 59929
rect 10355 59915 10407 59929
rect 10407 59915 10409 59929
rect 10353 59877 10355 59891
rect 10355 59877 10407 59891
rect 10407 59877 10409 59891
rect 10353 59865 10409 59877
rect 10353 59835 10355 59865
rect 10355 59835 10407 59865
rect 10407 59835 10409 59865
rect 27058 59066 27514 59522
rect 15411 57229 16507 57365
rect -377 56893 -321 56949
rect -297 56893 -241 56949
rect -217 56893 -161 56949
rect -137 56893 -81 56949
rect -57 56893 -1 56949
rect 23 56893 79 56949
rect 103 56893 159 56949
rect 41898 57449 42594 57585
rect 17618 57180 18794 57316
rect 43234 57162 43930 57171
rect 43234 57046 43256 57162
rect 43256 57046 43930 57162
rect 43234 57035 43930 57046
rect 16584 55639 17280 55775
rect 28024 55774 28800 55784
rect 28024 55658 28034 55774
rect 28034 55658 28790 55774
rect 28790 55658 28800 55774
rect 28024 55648 28800 55658
rect 13020 55242 13636 55378
rect 10150 53186 10152 53216
rect 10152 53186 10204 53216
rect 10204 53186 10206 53216
rect 10150 53174 10206 53186
rect 10150 53160 10152 53174
rect 10152 53160 10204 53174
rect 10204 53160 10206 53174
rect 10150 53122 10152 53136
rect 10152 53122 10204 53136
rect 10204 53122 10206 53136
rect 10150 53110 10206 53122
rect 10150 53080 10152 53110
rect 10152 53080 10204 53110
rect 10204 53080 10206 53110
rect -364 50128 172 50264
rect 9962 46451 9964 46481
rect 9964 46451 10016 46481
rect 10016 46451 10018 46481
rect 9962 46439 10018 46451
rect 9962 46425 9964 46439
rect 9964 46425 10016 46439
rect 10016 46425 10018 46439
rect 9962 46387 9964 46401
rect 9964 46387 10016 46401
rect 10016 46387 10018 46401
rect 9962 46375 10018 46387
rect 9962 46345 9964 46375
rect 9964 46345 10016 46375
rect 10016 46345 10018 46375
rect -378 43447 -322 43503
rect -298 43447 -242 43503
rect -218 43447 -162 43503
rect -138 43447 -82 43503
rect -58 43447 -2 43503
rect 22 43447 78 43503
rect 102 43447 158 43503
rect 9762 39738 9764 39768
rect 9764 39738 9816 39768
rect 9816 39738 9818 39768
rect 9762 39726 9818 39738
rect 9762 39712 9764 39726
rect 9764 39712 9816 39726
rect 9816 39712 9818 39726
rect 9762 39674 9764 39688
rect 9764 39674 9816 39688
rect 9816 39674 9818 39688
rect 9762 39662 9818 39674
rect 9762 39632 9764 39662
rect 9764 39632 9816 39662
rect 9816 39632 9818 39662
rect -377 36724 159 36860
rect 9539 32938 9541 32968
rect 9541 32938 9593 32968
rect 9593 32938 9595 32968
rect 9539 32926 9595 32938
rect 9539 32912 9541 32926
rect 9541 32912 9593 32926
rect 9593 32912 9595 32926
rect 9539 32874 9541 32888
rect 9541 32874 9593 32888
rect 9593 32874 9595 32888
rect 9539 32862 9595 32874
rect 9539 32832 9541 32862
rect 9541 32832 9593 32862
rect 9593 32832 9595 32862
rect -379 29941 157 30077
rect 8520 26010 8522 26040
rect 8522 26010 8574 26040
rect 8574 26010 8576 26040
rect 8520 25998 8576 26010
rect 8520 25984 8522 25998
rect 8522 25984 8574 25998
rect 8574 25984 8576 25998
rect 8520 25946 8522 25960
rect 8522 25946 8574 25960
rect 8574 25946 8576 25960
rect 8520 25934 8576 25946
rect 8520 25904 8522 25934
rect 8522 25904 8574 25934
rect 8574 25904 8576 25934
rect -364 23015 -308 23071
rect -284 23015 -228 23071
rect -204 23015 -148 23071
rect -124 23015 -68 23071
rect -44 23015 12 23071
rect 36 23015 92 23071
rect 116 23015 172 23071
rect 8724 19370 8780 19380
rect 8724 19324 8726 19370
rect 8726 19324 8778 19370
rect 8778 19324 8780 19370
rect 8724 19254 8726 19300
rect 8726 19254 8778 19300
rect 8778 19254 8780 19300
rect 8724 19244 8780 19254
rect -376 16281 -320 16337
rect -296 16281 -240 16337
rect -216 16281 -160 16337
rect -136 16281 -80 16337
rect -56 16281 0 16337
rect 24 16281 80 16337
rect 104 16281 160 16337
rect 8918 12557 8974 12567
rect 8918 12511 8920 12557
rect 8920 12511 8972 12557
rect 8972 12511 8974 12557
rect 8918 12441 8920 12487
rect 8920 12441 8972 12487
rect 8972 12441 8974 12487
rect 8918 12431 8974 12441
rect -374 9578 -318 9634
rect -294 9578 -238 9634
rect -214 9578 -158 9634
rect -134 9578 -78 9634
rect -54 9578 2 9634
rect 26 9578 82 9634
rect 106 9578 162 9634
rect 9120 5960 9176 5970
rect 9120 5914 9122 5960
rect 9122 5914 9174 5960
rect 9174 5914 9176 5960
rect 9120 5844 9122 5890
rect 9122 5844 9174 5890
rect 9174 5844 9176 5890
rect 9120 5834 9176 5844
rect -380 2844 156 2980
rect 9331 -863 9333 -833
rect 9333 -863 9385 -833
rect 9385 -863 9387 -833
rect 9331 -875 9387 -863
rect 9331 -889 9333 -875
rect 9333 -889 9385 -875
rect 9385 -889 9387 -875
rect 9331 -927 9333 -913
rect 9333 -927 9385 -913
rect 9385 -927 9387 -913
rect 9331 -939 9387 -927
rect 9331 -969 9333 -939
rect 9333 -969 9385 -939
rect 9385 -969 9387 -939
rect -377 -3950 159 -3814
rect 1809 -4644 1811 -4428
rect 1811 -4644 2183 -4428
rect 2183 -4644 2185 -4428
<< metal3 >>
rect 200 68131 66589 68178
rect 200 68122 64735 68131
rect 200 67666 36052 68122
rect 36348 67667 64735 68122
rect 64959 67667 66589 68131
rect 36348 67666 66589 67667
rect 200 67588 66589 67666
rect 33776 67410 34206 67436
rect 188 67373 66595 67410
rect 188 66917 33842 67373
rect 34138 67341 66595 67373
rect 34138 66917 65153 67341
rect 188 66877 65153 66917
rect 65377 66877 66595 67341
rect 188 66820 66595 66877
rect 26994 66588 27586 66616
rect 206 66548 66595 66588
rect 206 66485 27063 66548
rect 206 66181 15756 66485
rect 16220 66181 27063 66485
rect 206 66172 27063 66181
rect 27519 66526 66595 66548
rect 27519 66172 41828 66526
rect 206 66062 41828 66172
rect 42532 66473 66595 66526
rect 42532 66089 65696 66473
rect 65840 66089 66595 66473
rect 42532 66062 66595 66089
rect 206 65998 66595 66062
rect 196 65802 404 65814
rect 190 65735 66617 65802
rect 190 65271 18357 65735
rect 18901 65734 66617 65735
rect 18901 65271 43512 65734
rect 190 65270 43512 65271
rect 44216 65730 66617 65734
rect 44216 65270 66271 65730
rect 190 65266 66271 65270
rect 66495 65266 66617 65730
rect 190 65212 66617 65266
rect 29746 63435 31106 63474
rect 29746 63299 29796 63435
rect 31052 63299 31106 63435
rect 29746 63248 31106 63299
rect 30106 63244 30656 63248
rect 35992 62694 36416 62776
rect 35992 62477 36049 62694
rect 31245 62398 36049 62477
rect 36345 62398 36416 62694
rect 31245 62330 36416 62398
rect 31245 62319 36395 62330
rect 10320 59975 10452 60010
rect 10320 59911 10349 59975
rect 10413 59911 10452 59975
rect 10320 59895 10452 59911
rect 10320 59831 10349 59895
rect 10413 59831 10452 59895
rect 10320 59790 10452 59831
rect 26976 59522 27622 59608
rect 26976 59066 27058 59522
rect 27514 59211 27622 59522
rect 27514 59066 30915 59211
rect 26976 58990 30915 59066
rect 26985 58985 30915 58990
rect 41810 57589 42702 57628
rect 41810 57445 41894 57589
rect 42598 57445 42702 57589
rect 15380 57369 16564 57404
rect 41810 57382 42702 57445
rect 15380 57225 15407 57369
rect 16511 57225 16564 57369
rect 15380 57188 16564 57225
rect 17566 57320 18858 57362
rect 17566 57316 17654 57320
rect 18758 57316 18858 57320
rect 17566 57180 17618 57316
rect 18794 57180 18858 57316
rect 17566 57176 17654 57180
rect 18758 57176 18858 57180
rect 17566 57152 18858 57176
rect 43182 57175 43984 57204
rect 43182 57031 43230 57175
rect 43934 57031 43984 57175
rect 43182 57014 43984 57031
rect -400 56949 198 57004
rect -400 56893 -377 56949
rect -321 56893 -297 56949
rect -241 56893 -217 56949
rect -161 56893 -137 56949
rect -81 56893 -57 56949
rect -1 56893 23 56949
rect 79 56893 103 56949
rect 159 56893 198 56949
rect -400 56836 198 56893
rect 10804 55784 47572 55808
rect 10804 55778 28024 55784
rect 10804 55775 19038 55778
rect 10804 55639 16584 55775
rect 17280 55639 19038 55775
rect 10804 55634 19038 55639
rect 19742 55648 28024 55778
rect 28800 55648 47572 55784
rect 19742 55634 47572 55648
rect 10804 55602 47572 55634
rect 12984 55382 13674 55428
rect 12984 55238 13016 55382
rect 13640 55238 13674 55382
rect 12984 55206 13674 55238
rect 66196 53775 66590 53834
rect 66196 53576 66301 53775
rect 61178 53376 66301 53576
rect 10118 53220 10236 53256
rect 10118 53156 10146 53220
rect 10210 53156 10236 53220
rect 10118 53140 10236 53156
rect 10118 53076 10146 53140
rect 10210 53076 10236 53140
rect 10118 53038 10236 53076
rect 66196 53151 66301 53376
rect 66525 53151 66590 53775
rect 66196 53058 66590 53151
rect -400 50264 206 50276
rect -400 50128 -364 50264
rect 172 50128 206 50264
rect -400 50102 206 50128
rect 9912 46485 10050 46512
rect 9912 46421 9958 46485
rect 10022 46421 10050 46485
rect 9912 46405 10050 46421
rect 9912 46341 9958 46405
rect 10022 46341 10050 46405
rect 9912 46304 10050 46341
rect -402 43503 198 43554
rect -402 43447 -378 43503
rect -322 43447 -298 43503
rect -242 43447 -218 43503
rect -162 43447 -138 43503
rect -82 43447 -58 43503
rect -2 43447 22 43503
rect 78 43447 102 43503
rect 158 43447 198 43503
rect -402 43388 198 43447
rect 8484 40803 11003 40840
rect 8484 40739 10343 40803
rect 10407 40739 11003 40803
rect 8484 40723 11003 40739
rect 8484 40659 10343 40723
rect 10407 40659 11003 40723
rect 8484 40622 11003 40659
rect 8488 40428 11004 40462
rect 8488 40364 10149 40428
rect 10213 40364 11004 40428
rect 8488 40348 11004 40364
rect 8488 40284 10149 40348
rect 10213 40284 11004 40348
rect 8488 40244 11004 40284
rect 9728 39772 9854 39804
rect 9728 39708 9758 39772
rect 9822 39708 9854 39772
rect 9728 39692 9854 39708
rect 9728 39628 9758 39692
rect 9822 39628 9854 39692
rect 9728 39588 9854 39628
rect -402 36860 204 36870
rect -402 36724 -377 36860
rect 159 36724 204 36860
rect -402 36700 204 36724
rect 8490 35124 10990 35152
rect 8490 35060 9956 35124
rect 10020 35060 10990 35124
rect 8490 35044 10990 35060
rect 8490 34980 9956 35044
rect 10020 34980 10990 35044
rect 8490 34936 10990 34980
rect 8492 34758 11004 34770
rect 8488 34726 11124 34758
rect 8488 34662 9754 34726
rect 9818 34662 11124 34726
rect 8488 34646 11124 34662
rect 8488 34582 9754 34646
rect 9818 34582 11124 34646
rect 8488 34550 11124 34582
rect 9502 32972 9632 33008
rect 9502 32908 9535 32972
rect 9599 32908 9632 32972
rect 9502 32892 9632 32908
rect 9502 32828 9535 32892
rect 9599 32828 9632 32892
rect 9502 32790 9632 32828
rect -416 30077 206 30094
rect -416 29941 -379 30077
rect 157 29941 206 30077
rect -416 29922 206 29941
rect 8482 29398 11404 29430
rect 782 29371 956 29384
rect -414 29173 196 29200
rect -414 29029 -386 29173
rect 158 29029 196 29173
rect -414 28996 196 29029
rect 782 28907 797 29371
rect 941 28907 956 29371
rect 8482 29334 9533 29398
rect 9597 29334 11404 29398
rect 8482 29318 11404 29334
rect 8482 29254 9533 29318
rect 9597 29254 11404 29318
rect 8482 29216 11404 29254
rect 782 28894 956 28907
rect 8480 29030 11012 29036
rect 8480 29003 11026 29030
rect 8480 28939 8512 29003
rect 8576 28939 11026 29003
rect 8480 28923 11026 28939
rect 8480 28859 8512 28923
rect 8576 28859 11026 28923
rect 8480 28828 11026 28859
rect 8494 28822 11026 28828
rect -400 28748 586 28750
rect -408 28522 586 28748
rect -408 28520 210 28522
rect 8488 26044 8604 26070
rect 8488 25980 8516 26044
rect 8580 25980 8604 26044
rect 8488 25964 8604 25980
rect 8488 25900 8516 25964
rect 8580 25900 8604 25964
rect 8488 25864 8604 25900
rect 8490 23790 10858 23816
rect 8490 23726 8706 23790
rect 8770 23726 10858 23790
rect 8490 23710 10858 23726
rect 8490 23646 8706 23710
rect 8770 23646 10858 23710
rect 8490 23614 10858 23646
rect 8484 23400 10894 23430
rect 8484 23336 8920 23400
rect 8984 23336 10894 23400
rect 8484 23320 10894 23336
rect 8484 23256 8920 23320
rect 8984 23256 10894 23320
rect 8484 23224 10894 23256
rect -400 23071 198 23124
rect -400 23015 -364 23071
rect -308 23015 -284 23071
rect -228 23015 -204 23071
rect -148 23015 -124 23071
rect -68 23015 -44 23071
rect 12 23015 36 23071
rect 92 23015 116 23071
rect 172 23015 198 23071
rect -400 22950 198 23015
rect 8690 19384 8812 19406
rect 8690 19320 8720 19384
rect 8784 19320 8812 19384
rect 8690 19304 8812 19320
rect 8690 19240 8720 19304
rect 8784 19240 8812 19304
rect 8690 19210 8812 19240
rect 8482 18127 11328 18150
rect 8482 18063 9109 18127
rect 9173 18063 11328 18127
rect 8482 18047 11328 18063
rect 8482 17983 9109 18047
rect 9173 17983 11328 18047
rect 8482 17950 11328 17983
rect 8484 17686 12158 17710
rect 8484 17622 9331 17686
rect 9395 17622 12158 17686
rect 8484 17606 12158 17622
rect 8484 17542 9331 17606
rect 9395 17542 12158 17606
rect 8484 17510 12158 17542
rect -404 16337 196 16392
rect -404 16281 -376 16337
rect -320 16281 -296 16337
rect -240 16281 -216 16337
rect -160 16281 -136 16337
rect -80 16281 -56 16337
rect 0 16281 24 16337
rect 80 16281 104 16337
rect 160 16281 196 16337
rect -404 16224 196 16281
rect 8890 12571 9008 12598
rect 8890 12507 8914 12571
rect 8978 12507 9008 12571
rect 8890 12491 9008 12507
rect 8890 12427 8914 12491
rect 8978 12427 9008 12491
rect 8890 12394 9008 12427
rect -410 9634 200 9680
rect -410 9578 -374 9634
rect -318 9578 -294 9634
rect -238 9578 -214 9634
rect -158 9578 -134 9634
rect -78 9578 -54 9634
rect 2 9578 26 9634
rect 82 9578 106 9634
rect 162 9578 200 9634
rect -410 9510 200 9578
rect 9086 5974 9200 6002
rect 9086 5910 9116 5974
rect 9180 5910 9200 5974
rect 9086 5894 9200 5910
rect 9086 5830 9116 5894
rect 9180 5830 9200 5894
rect 9086 5798 9200 5830
rect 66220 5081 66574 5172
rect 66220 5020 66292 5081
rect 61363 4814 66292 5020
rect 66220 4697 66292 4814
rect 66516 5020 66574 5081
rect 66516 4814 66601 5020
rect 66516 4697 66574 4814
rect 66220 4612 66574 4697
rect -402 2980 196 2992
rect -402 2844 -380 2980
rect 156 2844 196 2980
rect -402 2816 196 2844
rect 9298 -829 9416 -786
rect 9298 -893 9327 -829
rect 9391 -893 9416 -829
rect 9298 -909 9416 -893
rect 9298 -973 9327 -909
rect 9391 -973 9416 -909
rect 9298 -1012 9416 -973
rect -404 -3814 200 -3794
rect -404 -3950 -377 -3814
rect 159 -3950 200 -3814
rect -404 -3968 200 -3950
rect 1750 -4424 2216 -4374
rect 1750 -4648 1805 -4424
rect 2189 -4648 2216 -4424
rect 1750 -4738 2216 -4648
rect 2482 -4474 3010 -4426
rect 2482 -4618 2540 -4474
rect 2924 -4618 3010 -4474
rect 2482 -4714 3010 -4618
rect 5458 -4443 6400 -4386
rect 5458 -4747 5520 -4443
rect 6304 -4747 6400 -4443
rect 5458 -4788 6400 -4747
rect -946 -5112 492 -5094
rect -946 -5139 66602 -5112
rect -946 -5174 64672 -5139
rect -946 -5398 2529 -5174
rect 2913 -5398 64672 -5174
rect -946 -5443 64672 -5398
rect 64976 -5443 66602 -5139
rect -946 -5488 66602 -5443
rect -946 -5504 492 -5488
rect -930 -5666 66618 -5664
rect -946 -5709 66618 -5666
rect -946 -5750 65142 -5709
rect -946 -5974 1802 -5750
rect 2186 -5974 65142 -5750
rect -946 -6013 65142 -5974
rect 65446 -6013 66618 -5709
rect -946 -6028 66618 -6013
rect -930 -6040 66618 -6028
rect -928 -6166 528 -6152
rect -930 -6199 66618 -6166
rect -930 -6423 5548 -6199
rect 6332 -6423 65632 -6199
rect -930 -6503 5628 -6423
rect 5932 -6503 65632 -6423
rect 65936 -6503 66618 -6199
rect -930 -6542 66618 -6503
rect -932 -6714 516 -6700
rect -938 -6790 66608 -6714
rect -938 -7014 66231 -6790
rect 66535 -7014 66608 -6790
rect -938 -7090 66608 -7014
<< via3 >>
rect 64735 67667 64959 68131
rect 65153 66877 65377 67341
rect 15756 66181 16220 66485
rect 41828 66062 42532 66526
rect 65696 66089 65840 66473
rect 18357 65271 18901 65735
rect 43512 65270 44216 65734
rect 66271 65266 66495 65730
rect 10349 59971 10413 59975
rect 10349 59915 10353 59971
rect 10353 59915 10409 59971
rect 10409 59915 10413 59971
rect 10349 59911 10413 59915
rect 10349 59891 10413 59895
rect 10349 59835 10353 59891
rect 10353 59835 10409 59891
rect 10409 59835 10413 59891
rect 10349 59831 10413 59835
rect 41894 57585 42598 57589
rect 41894 57449 41898 57585
rect 41898 57449 42594 57585
rect 42594 57449 42598 57585
rect 41894 57445 42598 57449
rect 15407 57365 16511 57369
rect 15407 57229 15411 57365
rect 15411 57229 16507 57365
rect 16507 57229 16511 57365
rect 15407 57225 16511 57229
rect 17654 57316 18758 57320
rect 17654 57180 18758 57316
rect 17654 57176 18758 57180
rect 43230 57171 43934 57175
rect 43230 57035 43234 57171
rect 43234 57035 43930 57171
rect 43930 57035 43934 57171
rect 43230 57031 43934 57035
rect 19038 55634 19742 55778
rect 13016 55378 13640 55382
rect 13016 55242 13020 55378
rect 13020 55242 13636 55378
rect 13636 55242 13640 55378
rect 13016 55238 13640 55242
rect 10146 53216 10210 53220
rect 10146 53160 10150 53216
rect 10150 53160 10206 53216
rect 10206 53160 10210 53216
rect 10146 53156 10210 53160
rect 10146 53136 10210 53140
rect 10146 53080 10150 53136
rect 10150 53080 10206 53136
rect 10206 53080 10210 53136
rect 10146 53076 10210 53080
rect 66301 53151 66525 53775
rect 9958 46481 10022 46485
rect 9958 46425 9962 46481
rect 9962 46425 10018 46481
rect 10018 46425 10022 46481
rect 9958 46421 10022 46425
rect 9958 46401 10022 46405
rect 9958 46345 9962 46401
rect 9962 46345 10018 46401
rect 10018 46345 10022 46401
rect 9958 46341 10022 46345
rect 10343 40739 10407 40803
rect 10343 40659 10407 40723
rect 10149 40364 10213 40428
rect 10149 40284 10213 40348
rect 9758 39768 9822 39772
rect 9758 39712 9762 39768
rect 9762 39712 9818 39768
rect 9818 39712 9822 39768
rect 9758 39708 9822 39712
rect 9758 39688 9822 39692
rect 9758 39632 9762 39688
rect 9762 39632 9818 39688
rect 9818 39632 9822 39688
rect 9758 39628 9822 39632
rect 9956 35060 10020 35124
rect 9956 34980 10020 35044
rect 9754 34662 9818 34726
rect 9754 34582 9818 34646
rect 9535 32968 9599 32972
rect 9535 32912 9539 32968
rect 9539 32912 9595 32968
rect 9595 32912 9599 32968
rect 9535 32908 9599 32912
rect 9535 32888 9599 32892
rect 9535 32832 9539 32888
rect 9539 32832 9595 32888
rect 9595 32832 9599 32888
rect 9535 32828 9599 32832
rect -386 29029 158 29173
rect 797 28907 941 29371
rect 9533 29334 9597 29398
rect 9533 29254 9597 29318
rect 8512 28939 8576 29003
rect 8512 28859 8576 28923
rect 8516 26040 8580 26044
rect 8516 25984 8520 26040
rect 8520 25984 8576 26040
rect 8576 25984 8580 26040
rect 8516 25980 8580 25984
rect 8516 25960 8580 25964
rect 8516 25904 8520 25960
rect 8520 25904 8576 25960
rect 8576 25904 8580 25960
rect 8516 25900 8580 25904
rect 8706 23726 8770 23790
rect 8706 23646 8770 23710
rect 8920 23336 8984 23400
rect 8920 23256 8984 23320
rect 8720 19380 8784 19384
rect 8720 19324 8724 19380
rect 8724 19324 8780 19380
rect 8780 19324 8784 19380
rect 8720 19320 8784 19324
rect 8720 19300 8784 19304
rect 8720 19244 8724 19300
rect 8724 19244 8780 19300
rect 8780 19244 8784 19300
rect 8720 19240 8784 19244
rect 9109 18063 9173 18127
rect 9109 17983 9173 18047
rect 9331 17622 9395 17686
rect 9331 17542 9395 17606
rect 8914 12567 8978 12571
rect 8914 12511 8918 12567
rect 8918 12511 8974 12567
rect 8974 12511 8978 12567
rect 8914 12507 8978 12511
rect 8914 12487 8978 12491
rect 8914 12431 8918 12487
rect 8918 12431 8974 12487
rect 8974 12431 8978 12487
rect 8914 12427 8978 12431
rect 9116 5970 9180 5974
rect 9116 5914 9120 5970
rect 9120 5914 9176 5970
rect 9176 5914 9180 5970
rect 9116 5910 9180 5914
rect 9116 5890 9180 5894
rect 9116 5834 9120 5890
rect 9120 5834 9176 5890
rect 9176 5834 9180 5890
rect 9116 5830 9180 5834
rect 66292 4697 66516 5081
rect 9327 -833 9391 -829
rect 9327 -889 9331 -833
rect 9331 -889 9387 -833
rect 9387 -889 9391 -833
rect 9327 -893 9391 -889
rect 9327 -913 9391 -909
rect 9327 -969 9331 -913
rect 9331 -969 9387 -913
rect 9387 -969 9391 -913
rect 9327 -973 9391 -969
rect 1805 -4428 2189 -4424
rect 1805 -4644 1809 -4428
rect 1809 -4644 2185 -4428
rect 2185 -4644 2189 -4428
rect 1805 -4648 2189 -4644
rect 2540 -4618 2924 -4474
rect 5520 -4747 6304 -4443
rect 2529 -5398 2913 -5174
rect 64672 -5443 64976 -5139
rect 1802 -5974 2186 -5750
rect 65142 -6013 65446 -5709
rect 5548 -6423 6332 -6199
rect 5628 -6503 5932 -6423
rect 65632 -6503 65936 -6199
rect 66231 -7014 66535 -6790
<< metal4 >>
rect 15708 66485 16282 68183
rect 15708 66181 15756 66485
rect 16220 66181 16282 66485
rect 758 29371 982 29426
rect 758 29204 797 29371
rect -406 29173 797 29204
rect -406 29029 -386 29173
rect 158 29029 797 29173
rect -406 28996 797 29029
rect 758 28907 797 28996
rect 941 28907 982 29371
rect 758 28842 982 28907
rect 8488 29003 8608 62116
rect 8488 28939 8512 29003
rect 8576 28939 8608 29003
rect 8488 28923 8608 28939
rect 8488 28859 8512 28923
rect 8576 28859 8608 28923
rect 8488 26044 8608 28859
rect 8488 25980 8516 26044
rect 8580 25980 8608 26044
rect 8488 25964 8608 25980
rect 8488 25900 8516 25964
rect 8580 25900 8608 25964
rect 1750 -4424 2232 -4374
rect 1750 -4648 1805 -4424
rect 2189 -4648 2232 -4424
rect 1750 -4738 2232 -4648
rect 1756 -5750 2232 -4738
rect 2476 -4474 2998 -4426
rect 2476 -4618 2540 -4474
rect 2924 -4618 2998 -4474
rect 2476 -5174 2998 -4618
rect 2476 -5398 2529 -5174
rect 2913 -5398 2998 -5174
rect 2476 -5488 2998 -5398
rect 5458 -4443 6406 -4386
rect 5458 -4747 5520 -4443
rect 6304 -4747 6406 -4443
rect 8488 -4626 8608 25900
rect 8690 23790 8810 62116
rect 8690 23726 8706 23790
rect 8770 23726 8810 23790
rect 8690 23710 8810 23726
rect 8690 23646 8706 23710
rect 8770 23646 8810 23710
rect 8690 19384 8810 23646
rect 8690 19320 8720 19384
rect 8784 19320 8810 19384
rect 8690 19304 8810 19320
rect 8690 19240 8720 19304
rect 8784 19240 8810 19304
rect 8690 -4626 8810 19240
rect 8892 23400 9012 62116
rect 8892 23336 8920 23400
rect 8984 23336 9012 23400
rect 8892 23320 9012 23336
rect 8892 23256 8920 23320
rect 8984 23256 9012 23320
rect 8892 12598 9012 23256
rect 8890 12571 9012 12598
rect 8890 12507 8914 12571
rect 8978 12507 9012 12571
rect 8890 12491 9012 12507
rect 8890 12427 8914 12491
rect 8978 12427 9012 12491
rect 8890 12394 9012 12427
rect 8892 -4626 9012 12394
rect 9086 18127 9206 62116
rect 9086 18063 9109 18127
rect 9173 18063 9206 18127
rect 9086 18047 9206 18063
rect 9086 17983 9109 18047
rect 9173 17983 9206 18047
rect 9086 5974 9206 17983
rect 9086 5910 9116 5974
rect 9180 5910 9206 5974
rect 9086 5894 9206 5910
rect 9086 5830 9116 5894
rect 9180 5830 9206 5894
rect 9086 -4626 9206 5830
rect 9306 17686 9426 62116
rect 9306 17622 9331 17686
rect 9395 17622 9426 17686
rect 9306 17606 9426 17622
rect 9306 17542 9331 17606
rect 9395 17542 9426 17606
rect 9306 -786 9426 17542
rect 9298 -829 9426 -786
rect 9298 -893 9327 -829
rect 9391 -893 9426 -829
rect 9298 -909 9426 -893
rect 9298 -973 9327 -909
rect 9391 -973 9426 -909
rect 9298 -1012 9426 -973
rect 9306 -4626 9426 -1012
rect 9506 32972 9626 62116
rect 9506 32908 9535 32972
rect 9599 32908 9626 32972
rect 9506 32892 9626 32908
rect 9506 32828 9535 32892
rect 9599 32828 9626 32892
rect 9506 29398 9626 32828
rect 9506 29334 9533 29398
rect 9597 29334 9626 29398
rect 9506 29318 9626 29334
rect 9506 29254 9533 29318
rect 9597 29254 9626 29318
rect 9506 -4626 9626 29254
rect 9730 39772 9850 62116
rect 9730 39708 9758 39772
rect 9822 39708 9850 39772
rect 9730 39692 9850 39708
rect 9730 39628 9758 39692
rect 9822 39628 9850 39692
rect 9730 34726 9850 39628
rect 9730 34662 9754 34726
rect 9818 34662 9850 34726
rect 9730 34646 9850 34662
rect 9730 34582 9754 34646
rect 9818 34582 9850 34646
rect 9730 -4626 9850 34582
rect 9926 46485 10046 62116
rect 9926 46421 9958 46485
rect 10022 46421 10046 46485
rect 9926 46405 10046 46421
rect 9926 46341 9958 46405
rect 10022 46341 10046 46405
rect 9926 35124 10046 46341
rect 9926 35060 9956 35124
rect 10020 35060 10046 35124
rect 9926 35044 10046 35060
rect 9926 34980 9956 35044
rect 10020 34980 10046 35044
rect 9926 -4626 10046 34980
rect 10120 53220 10240 62116
rect 10120 53156 10146 53220
rect 10210 53156 10240 53220
rect 10120 53140 10240 53156
rect 10120 53076 10146 53140
rect 10210 53076 10240 53140
rect 10120 40428 10240 53076
rect 10120 40364 10149 40428
rect 10213 40364 10240 40428
rect 10120 40348 10240 40364
rect 10120 40284 10149 40348
rect 10213 40284 10240 40348
rect 10120 -4626 10240 40284
rect 10320 59975 10440 62116
rect 10320 59911 10349 59975
rect 10413 59911 10440 59975
rect 10320 59895 10440 59911
rect 10320 59831 10349 59895
rect 10413 59831 10440 59895
rect 10320 40803 10440 59831
rect 15708 57404 16282 66181
rect 18314 65735 18986 68198
rect 18314 65271 18357 65735
rect 18901 65271 18986 65735
rect 15380 57369 16564 57404
rect 18314 57372 18986 65271
rect 41786 66526 42584 68183
rect 41786 66062 41828 66526
rect 42532 66062 42584 66526
rect 41786 57874 42584 66062
rect 43390 65734 44270 68184
rect 43390 65270 43512 65734
rect 44216 65270 44270 65734
rect 41786 57792 42588 57874
rect 41794 57628 42588 57792
rect 41794 57589 42702 57628
rect 41794 57445 41894 57589
rect 42598 57445 42702 57589
rect 41794 57386 42702 57445
rect 41810 57382 42702 57386
rect 15380 57225 15407 57369
rect 16511 57225 16564 57369
rect 15380 57188 16564 57225
rect 17564 57320 18986 57372
rect 17564 57176 17654 57320
rect 18758 57176 18986 57320
rect 43390 57204 44270 65270
rect 17564 57134 18986 57176
rect 43182 57175 44270 57204
rect 43182 57031 43230 57175
rect 43934 57031 44270 57175
rect 43182 57022 44270 57031
rect 64642 68131 65018 68240
rect 64642 67667 64735 68131
rect 64959 67667 65018 68131
rect 43182 57014 43984 57022
rect 19244 55804 19448 55806
rect 18974 55778 19768 55804
rect 18974 55634 19038 55778
rect 19742 55634 19768 55778
rect 18974 55596 19768 55634
rect 12988 55382 13676 55408
rect 12988 55238 13016 55382
rect 13640 55238 13676 55382
rect 12988 55208 13676 55238
rect 13250 52206 13454 55208
rect 19244 51418 19448 55596
rect 10320 40739 10343 40803
rect 10407 40739 10440 40803
rect 10320 40723 10440 40739
rect 10320 40659 10343 40723
rect 10407 40659 10440 40723
rect 10320 -4626 10440 40659
rect 1756 -5974 1802 -5750
rect 2186 -5974 2232 -5750
rect 1756 -6042 2232 -5974
rect 5458 -6199 6406 -4747
rect 64642 -5084 65018 67667
rect 65112 67341 65488 68240
rect 65112 66877 65153 67341
rect 65377 66877 65488 67341
rect 64630 -5139 65030 -5084
rect 64630 -5443 64672 -5139
rect 64976 -5443 65030 -5139
rect 64630 -5484 65030 -5443
rect 5458 -6423 5548 -6199
rect 6332 -6423 6406 -6199
rect 5458 -6503 5628 -6423
rect 5932 -6503 6406 -6423
rect 5458 -6594 6406 -6503
rect 64642 -7084 65018 -5484
rect 65112 -5709 65488 66877
rect 65112 -6013 65142 -5709
rect 65446 -6013 65488 -5709
rect 65112 -7090 65488 -6013
rect 65592 66473 65968 68240
rect 65592 66089 65696 66473
rect 65840 66089 65968 66473
rect 65592 -6199 65968 66089
rect 65592 -6503 65632 -6199
rect 65936 -6503 65968 -6199
rect 65592 -7090 65968 -6503
rect 66208 65730 66584 68202
rect 66208 65266 66271 65730
rect 66495 65266 66584 65730
rect 66208 53775 66584 65266
rect 66208 53151 66301 53775
rect 66525 53151 66584 53775
rect 66208 5081 66584 53151
rect 66208 4697 66292 5081
rect 66516 4697 66584 5081
rect 66208 -6790 66584 4697
rect 66208 -7014 66231 -6790
rect 66535 -7014 66584 -6790
rect 66208 -7090 66584 -7014
use capbank_8b8  capbank_8b8_0
timestamp 1699926577
transform 1 0 13952 0 1 24020
box -3422 -20118 50401 30484
use EF_AMUX21_ARRAY  EF_AMUX21_ARRAY_0
timestamp 1699926577
transform 0 1 1180 -1 0 14388
box -49267 -1504 20268 7804
use EF_BUF3V3  EF_BUF3V3_0
timestamp 1699926577
transform 0 -1 17605 1 0 61545
box -4547 -3901 2817 6641
use EF_BUF3V3  EF_BUF3V3_1
timestamp 1699926577
transform 0 -1 43613 1 0 61759
box -4547 -3901 2817 6641
use EF_SW_RST  EF_SW_RST_1
timestamp 1699926577
transform 1 0 32340 0 -1 63067
box -5689 -398 2820 6071
<< labels >>
flabel metal3 s -946 -5504 492 -5094 0 FreeSans 3601 0 0 0 DVDD
port 1 nsew
flabel metal3 s -946 -6028 510 -5666 0 FreeSans 3601 0 0 0 DVSS
port 2 nsew
flabel metal3 s -928 -6514 528 -6152 0 FreeSans 3601 0 0 0 VDD
port 3 nsew
flabel metal3 s -932 -7074 516 -6700 0 FreeSans 12631 0 0 0 VSS
port 4 nsew
flabel metal2 s 21622 68364 21822 68924 0 FreeSans 10105 0 0 0 EN
port 5 nsew
flabel metal2 s 17200 68318 17432 68986 0 FreeSans 8083 0 0 0 OUT
port 6 nsew
flabel metal2 s 30190 68212 30412 68814 0 FreeSans 4139 0 0 0 RST
port 7 nsew
flabel metal3 s -414 28996 196 29200 0 FreeSans 3476 0 0 0 VH
port 8 nsew
flabel metal3 s -408 28520 210 28748 0 FreeSans 3476 0 0 0 VL
port 9 nsew
flabel metal3 s -416 29922 206 30094 0 FreeSans 3476 0 0 0 SELD5
port 10 nsew
flabel metal3 s -400 22950 198 23124 0 FreeSans 1736 0 0 0 SELD0
port 11 nsew
flabel metal3 s -404 16224 196 16392 0 FreeSans 1736 0 0 0 SELD1
port 12 nsew
flabel metal3 s -410 9510 200 9680 0 FreeSans 1736 0 0 0 SELD2
port 13 nsew
flabel metal3 s -402 2816 196 2992 0 FreeSans 1736 0 0 0 SELD3
port 14 nsew
flabel metal3 s -404 -3968 200 -3794 0 FreeSans 1736 0 0 0 SELD4
port 15 nsew
flabel metal3 s -400 56836 198 57004 0 FreeSans 1736 0 0 0 SELD9
port 16 nsew
flabel metal3 s -400 50102 206 50276 0 FreeSans 1736 0 0 0 SELD8
port 17 nsew
flabel metal3 s -402 43388 198 43554 0 FreeSans 1736 0 0 0 SELD7
port 18 nsew
flabel metal3 s -402 36700 204 36870 0 FreeSans 1736 0 0 0 SELD6
port 19 nsew
<< end >>
