magic
tech sky130A
magscale 1 2
timestamp 1693827120
<< metal3 >>
rect -650 552 731 600
rect -650 488 647 552
rect 711 488 731 552
rect -650 472 731 488
rect -650 408 647 472
rect 711 408 731 472
rect -650 392 731 408
rect -650 328 647 392
rect 711 328 731 392
rect -650 312 731 328
rect -650 248 647 312
rect 711 248 731 312
rect -650 232 731 248
rect -650 168 647 232
rect 711 168 731 232
rect -650 152 731 168
rect -650 88 647 152
rect 711 88 731 152
rect -650 72 731 88
rect -650 8 647 72
rect 711 8 731 72
rect -650 -8 731 8
rect -650 -72 647 -8
rect 711 -72 731 -8
rect -650 -88 731 -72
rect -650 -152 647 -88
rect 711 -152 731 -88
rect -650 -168 731 -152
rect -650 -232 647 -168
rect 711 -232 731 -168
rect -650 -248 731 -232
rect -650 -312 647 -248
rect 711 -312 731 -248
rect -650 -328 731 -312
rect -650 -392 647 -328
rect 711 -392 731 -328
rect -650 -408 731 -392
rect -650 -472 647 -408
rect 711 -472 731 -408
rect -650 -488 731 -472
rect -650 -552 647 -488
rect 711 -552 731 -488
rect -650 -600 731 -552
<< via3 >>
rect 647 488 711 552
rect 647 408 711 472
rect 647 328 711 392
rect 647 248 711 312
rect 647 168 711 232
rect 647 88 711 152
rect 647 8 711 72
rect 647 -72 711 -8
rect 647 -152 711 -88
rect 647 -232 711 -168
rect 647 -312 711 -248
rect 647 -392 711 -328
rect 647 -472 711 -408
rect 647 -552 711 -488
<< mimcap >>
rect -550 432 450 500
rect -550 -432 -482 432
rect 382 -432 450 432
rect -550 -500 450 -432
<< mimcapcontact >>
rect -482 -432 382 432
<< metal4 >>
rect 631 552 727 701
rect 631 488 647 552
rect 711 488 727 552
rect 631 472 727 488
rect -511 432 411 461
rect -511 -432 -482 432
rect 382 -432 411 432
rect -511 -461 411 -432
rect 631 408 647 472
rect 711 408 727 472
rect 631 392 727 408
rect 631 328 647 392
rect 711 328 727 392
rect 631 312 727 328
rect 631 248 647 312
rect 711 248 727 312
rect 631 232 727 248
rect 631 168 647 232
rect 711 168 727 232
rect 631 152 727 168
rect 631 88 647 152
rect 711 88 727 152
rect 631 72 727 88
rect 631 8 647 72
rect 711 8 727 72
rect 631 -8 727 8
rect 631 -72 647 -8
rect 711 -72 727 -8
rect 631 -88 727 -72
rect 631 -152 647 -88
rect 711 -152 727 -88
rect 631 -168 727 -152
rect 631 -232 647 -168
rect 711 -232 727 -168
rect 631 -248 727 -232
rect 631 -312 647 -248
rect 711 -312 727 -248
rect 631 -328 727 -312
rect 631 -392 647 -328
rect 711 -392 727 -328
rect 631 -408 727 -392
rect 631 -472 647 -408
rect 711 -472 727 -408
rect 631 -488 727 -472
rect 631 -552 647 -488
rect 711 -552 727 -488
rect 631 -588 727 -552
<< properties >>
string FIXED_BBOX -650 -600 550 600
<< end >>
