VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO EF_ADCS1008NC
  CLASS BLOCK ;
  FOREIGN EF_ADCS1008NC ;
  ORIGIN 0.000 0.000 ;
  SIZE 348.430 BY 531.590 ;
  PIN B[0]
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 179.120 500.640 180.660 500.940 ;
    END
  END B[0]
  PIN B[1]
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 179.110 499.950 180.650 500.250 ;
    END
  END B[1]
  PIN B[2]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 179.130 499.280 180.670 499.580 ;
    END
  END B[2]
  PIN VIN[0]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 144.370 530.050 144.825 531.540 ;
    END
  END VIN[0]
  PIN VIN[1]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 127.150 530.050 127.630 531.560 ;
    END
  END VIN[1]
  PIN VIN[2]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 110.630 530.070 111.110 531.580 ;
    END
  END VIN[2]
  PIN VIN[3]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 93.750 530.090 94.210 531.570 ;
    END
  END VIN[3]
  PIN VIN[4]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 77.200 530.060 77.660 531.540 ;
    END
  END VIN[4]
  PIN VIN[5]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 60.680 530.070 61.140 531.550 ;
    END
  END VIN[5]
  PIN VIN[6]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 43.690 530.070 44.150 531.550 ;
    END
  END VIN[6]
  PIN VIN[7]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 26.700 530.090 27.160 531.570 ;
    END
  END VIN[7]
  PIN HOLD
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT 10.430 447.815 11.430 448.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.570 447.830 7.720 448.840 ;
    END
  END HOLD
  PIN CMP
    ANTENNADIFFAREA 0.492900 ;
    PORT
      LAYER met3 ;
        RECT 178.550 424.110 180.620 425.100 ;
    END
  END CMP
  PIN DATA[9]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 10.580 333.580 16.340 334.460 ;
    END
  END DATA[9]
  PIN DATA[8]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 10.600 299.950 16.360 300.830 ;
    END
  END DATA[8]
  PIN DATA[7]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 10.560 266.370 16.320 267.250 ;
    END
  END DATA[7]
  PIN DATA[6]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 10.620 232.900 16.380 233.780 ;
    END
  END DATA[6]
  PIN DATA[5]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 10.640 199.050 16.400 199.930 ;
    END
  END DATA[5]
  PIN DATA[0]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 10.580 164.120 16.340 165.000 ;
    END
  END DATA[0]
  PIN DATA[1]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 10.620 130.590 16.380 131.470 ;
    END
  END DATA[1]
  PIN DATA[2]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 10.600 96.990 16.360 97.870 ;
    END
  END DATA[2]
  PIN DATA[3]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 10.560 63.480 16.320 64.360 ;
    END
  END DATA[3]
  PIN DATA[4]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 10.580 29.590 16.340 30.470 ;
    END
  END DATA[4]
  PIN VH
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met3 ;
        RECT 10.580 194.490 16.340 195.370 ;
    END
  END VH
  PIN VL
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met3 ;
        RECT 10.530 192.160 16.290 193.040 ;
    END
  END VL
  PIN RST
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER met3 ;
        RECT 8.580 391.130 12.680 392.140 ;
    END
  END RST
  PIN DVDD
    ANTENNAGATEAREA 47.261497 ;
    ANTENNADIFFAREA 93.596451 ;
    PORT
      LAYER met3 ;
        RECT 10.620 21.890 17.810 23.880 ;
    END
  END DVDD
  PIN DVSS
    ANTENNAGATEAREA 74.759102 ;
    ANTENNADIFFAREA 1023.766663 ;
    PORT
      LAYER met3 ;
        RECT 10.590 19.220 17.780 21.210 ;
    END
  END DVSS
  PIN VSS
    ANTENNAGATEAREA 130.500000 ;
    ANTENNADIFFAREA 621.362671 ;
    PORT
      LAYER met3 ;
        RECT 10.580 14.000 17.990 15.900 ;
    END
  END VSS
  PIN VDD
    ANTENNAGATEAREA 100.000000 ;
    ANTENNADIFFAREA 2509.495605 ;
    PORT
      LAYER met3 ;
        RECT 10.700 16.760 18.000 18.700 ;
    END
  END VDD
  PIN EN
    ANTENNAGATEAREA 1.752000 ;
    ANTENNADIFFAREA 1.080000 ;
    PORT
      LAYER met3 ;
        RECT 4.570 426.600 7.360 427.530 ;
    END
  END EN
  OBS
      LAYER li1 ;
        RECT 11.795 28.040 252.480 521.355 ;
      LAYER met1 ;
        RECT 4.615 449.095 253.175 521.560 ;
        RECT 4.615 447.535 10.150 449.095 ;
        RECT 11.710 447.535 253.175 449.095 ;
        RECT 4.615 25.725 253.175 447.535 ;
      LAYER met2 ;
        RECT 4.570 529.810 26.420 531.590 ;
        RECT 27.440 529.810 43.410 531.590 ;
        RECT 4.570 529.790 43.410 529.810 ;
        RECT 44.430 529.790 60.400 531.590 ;
        RECT 61.420 529.790 76.920 531.590 ;
        RECT 4.570 529.780 76.920 529.790 ;
        RECT 77.940 529.810 93.470 531.590 ;
        RECT 94.490 529.810 110.350 531.590 ;
        RECT 77.940 529.790 110.350 529.810 ;
        RECT 111.390 529.790 126.870 531.590 ;
        RECT 77.940 529.780 126.870 529.790 ;
        RECT 4.570 529.770 126.870 529.780 ;
        RECT 127.910 529.770 144.090 531.590 ;
        RECT 145.105 529.770 250.860 531.590 ;
        RECT 4.570 25.725 250.860 529.770 ;
      LAYER met3 ;
        RECT 4.560 501.340 348.430 529.560 ;
        RECT 4.560 500.650 178.720 501.340 ;
        RECT 4.560 499.550 178.710 500.650 ;
        RECT 181.060 500.240 348.430 501.340 ;
        RECT 181.050 499.980 348.430 500.240 ;
        RECT 4.560 498.880 178.730 499.550 ;
        RECT 181.070 498.880 348.430 499.980 ;
        RECT 4.560 449.240 348.430 498.880 ;
        RECT 8.120 447.430 348.430 449.240 ;
        RECT 4.560 427.930 348.430 447.430 ;
        RECT 7.760 426.200 348.430 427.930 ;
        RECT 4.560 425.500 348.430 426.200 ;
        RECT 4.560 423.710 178.150 425.500 ;
        RECT 181.020 423.710 348.430 425.500 ;
        RECT 4.560 392.540 348.430 423.710 ;
        RECT 4.560 390.730 8.180 392.540 ;
        RECT 13.080 390.730 348.430 392.540 ;
        RECT 4.560 334.860 348.430 390.730 ;
        RECT 4.560 333.180 10.180 334.860 ;
        RECT 16.740 333.180 348.430 334.860 ;
        RECT 4.560 301.230 348.430 333.180 ;
        RECT 4.560 299.550 10.200 301.230 ;
        RECT 16.760 299.550 348.430 301.230 ;
        RECT 4.560 267.650 348.430 299.550 ;
        RECT 4.560 265.970 10.160 267.650 ;
        RECT 16.720 265.970 348.430 267.650 ;
        RECT 4.560 234.180 348.430 265.970 ;
        RECT 4.560 232.500 10.220 234.180 ;
        RECT 16.780 232.500 348.430 234.180 ;
        RECT 4.560 200.330 348.430 232.500 ;
        RECT 4.560 198.650 10.240 200.330 ;
        RECT 16.800 198.650 348.430 200.330 ;
        RECT 4.560 195.770 348.430 198.650 ;
        RECT 4.560 194.090 10.180 195.770 ;
        RECT 16.740 194.090 348.430 195.770 ;
        RECT 4.560 193.440 348.430 194.090 ;
        RECT 4.560 191.760 10.130 193.440 ;
        RECT 16.690 191.760 348.430 193.440 ;
        RECT 4.560 165.400 348.430 191.760 ;
        RECT 4.560 163.720 10.180 165.400 ;
        RECT 16.740 163.720 348.430 165.400 ;
        RECT 4.560 131.870 348.430 163.720 ;
        RECT 4.560 130.190 10.220 131.870 ;
        RECT 16.780 130.190 348.430 131.870 ;
        RECT 4.560 98.270 348.430 130.190 ;
        RECT 4.560 96.590 10.200 98.270 ;
        RECT 16.760 96.590 348.430 98.270 ;
        RECT 4.560 64.760 348.430 96.590 ;
        RECT 4.560 63.080 10.160 64.760 ;
        RECT 16.720 63.080 348.430 64.760 ;
        RECT 4.560 30.870 348.430 63.080 ;
        RECT 4.560 29.190 10.180 30.870 ;
        RECT 16.740 29.190 348.430 30.870 ;
        RECT 4.560 24.280 348.430 29.190 ;
        RECT 4.560 21.610 10.220 24.280 ;
        RECT 4.560 18.820 10.190 21.610 ;
        RECT 18.210 21.490 348.430 24.280 ;
        RECT 18.180 19.100 348.430 21.490 ;
        RECT 4.560 16.360 10.300 18.820 ;
        RECT 18.400 16.360 348.430 19.100 ;
        RECT 4.560 16.300 348.430 16.360 ;
        RECT 4.560 13.965 10.180 16.300 ;
        RECT 18.390 13.965 348.430 16.300 ;
      LAYER met4 ;
        RECT 8.440 13.965 348.260 529.560 ;
      LAYER met5 ;
        RECT 21.505 398.445 175.535 520.875 ;
  END
END EF_ADCS1008NC
END LIBRARY

