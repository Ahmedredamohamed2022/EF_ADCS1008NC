magic
tech sky130A
magscale 1 2
timestamp 1699926577
<< nwell >>
rect -387 -362 387 362
<< mvpmos >>
rect -129 -64 -29 136
rect 29 -64 129 136
<< mvpdiff >>
rect -187 121 -129 136
rect -187 87 -175 121
rect -141 87 -129 121
rect -187 53 -129 87
rect -187 19 -175 53
rect -141 19 -129 53
rect -187 -15 -129 19
rect -187 -49 -175 -15
rect -141 -49 -129 -15
rect -187 -64 -129 -49
rect -29 121 29 136
rect -29 87 -17 121
rect 17 87 29 121
rect -29 53 29 87
rect -29 19 -17 53
rect 17 19 29 53
rect -29 -15 29 19
rect -29 -49 -17 -15
rect 17 -49 29 -15
rect -29 -64 29 -49
rect 129 121 187 136
rect 129 87 141 121
rect 175 87 187 121
rect 129 53 187 87
rect 129 19 141 53
rect 175 19 187 53
rect 129 -15 187 19
rect 129 -49 141 -15
rect 175 -49 187 -15
rect 129 -64 187 -49
<< mvpdiffc >>
rect -175 87 -141 121
rect -175 19 -141 53
rect -175 -49 -141 -15
rect -17 87 17 121
rect -17 19 17 53
rect -17 -49 17 -15
rect 141 87 175 121
rect 141 19 175 53
rect 141 -49 175 -15
<< mvnsubdiff >>
rect -321 284 321 296
rect -321 250 -187 284
rect -153 250 -119 284
rect -85 250 -51 284
rect -17 250 17 284
rect 51 250 85 284
rect 119 250 153 284
rect 187 250 321 284
rect -321 238 321 250
rect -321 187 -263 238
rect -321 153 -309 187
rect -275 153 -263 187
rect 263 187 321 238
rect -321 119 -263 153
rect 263 153 275 187
rect 309 153 321 187
rect -321 85 -309 119
rect -275 85 -263 119
rect -321 51 -263 85
rect -321 17 -309 51
rect -275 17 -263 51
rect -321 -17 -263 17
rect -321 -51 -309 -17
rect -275 -51 -263 -17
rect -321 -85 -263 -51
rect 263 119 321 153
rect 263 85 275 119
rect 309 85 321 119
rect 263 51 321 85
rect 263 17 275 51
rect 309 17 321 51
rect 263 -17 321 17
rect 263 -51 275 -17
rect 309 -51 321 -17
rect -321 -119 -309 -85
rect -275 -119 -263 -85
rect -321 -153 -263 -119
rect -321 -187 -309 -153
rect -275 -187 -263 -153
rect 263 -85 321 -51
rect 263 -119 275 -85
rect 309 -119 321 -85
rect 263 -153 321 -119
rect -321 -238 -263 -187
rect 263 -187 275 -153
rect 309 -187 321 -153
rect 263 -238 321 -187
rect -321 -250 321 -238
rect -321 -284 -187 -250
rect -153 -284 -119 -250
rect -85 -284 -51 -250
rect -17 -284 17 -250
rect 51 -284 85 -250
rect 119 -284 153 -250
rect 187 -284 321 -250
rect -321 -296 321 -284
<< mvnsubdiffcont >>
rect -187 250 -153 284
rect -119 250 -85 284
rect -51 250 -17 284
rect 17 250 51 284
rect 85 250 119 284
rect 153 250 187 284
rect -309 153 -275 187
rect 275 153 309 187
rect -309 85 -275 119
rect -309 17 -275 51
rect -309 -51 -275 -17
rect 275 85 309 119
rect 275 17 309 51
rect 275 -51 309 -17
rect -309 -119 -275 -85
rect -309 -187 -275 -153
rect 275 -119 309 -85
rect 275 -187 309 -153
rect -187 -284 -153 -250
rect -119 -284 -85 -250
rect -51 -284 -17 -250
rect 17 -284 51 -250
rect 85 -284 119 -250
rect 153 -284 187 -250
<< poly >>
rect -129 136 -29 162
rect 29 136 129 162
rect -129 -111 -29 -64
rect -129 -145 -96 -111
rect -62 -145 -29 -111
rect -129 -161 -29 -145
rect 29 -111 129 -64
rect 29 -145 62 -111
rect 96 -145 129 -111
rect 29 -161 129 -145
<< polycont >>
rect -96 -145 -62 -111
rect 62 -145 96 -111
<< locali >>
rect -309 250 -187 284
rect -153 250 -119 284
rect -85 250 -51 284
rect -17 250 17 284
rect 51 250 85 284
rect 119 250 153 284
rect 187 250 309 284
rect -309 187 -275 250
rect -309 119 -275 153
rect 275 187 309 250
rect -309 51 -275 85
rect -309 -17 -275 17
rect -309 -85 -275 -51
rect -175 121 -141 140
rect -175 53 -141 55
rect -175 17 -141 19
rect -175 -68 -141 -49
rect -17 121 17 140
rect -17 53 17 55
rect -17 17 17 19
rect -17 -68 17 -49
rect 141 121 175 140
rect 141 53 175 55
rect 141 17 175 19
rect 141 -68 175 -49
rect 275 119 309 153
rect 275 51 309 85
rect 275 -17 309 17
rect 275 -85 309 -51
rect -309 -153 -275 -119
rect -129 -145 -96 -111
rect -62 -145 -29 -111
rect 29 -145 62 -111
rect 96 -145 129 -111
rect -309 -250 -275 -187
rect 275 -153 309 -119
rect 275 -250 309 -187
rect -309 -284 -187 -250
rect -153 -284 -119 -250
rect -85 -284 -51 -250
rect -17 -284 17 -250
rect 51 -284 85 -250
rect 119 -284 153 -250
rect 187 -284 309 -250
<< viali >>
rect -175 87 -141 89
rect -175 55 -141 87
rect -175 -15 -141 17
rect -175 -17 -141 -15
rect -17 87 17 89
rect -17 55 17 87
rect -17 -15 17 17
rect -17 -17 17 -15
rect 141 87 175 89
rect 141 55 175 87
rect 141 -15 175 17
rect 141 -17 175 -15
rect -96 -145 -62 -111
rect 62 -145 96 -111
<< metal1 >>
rect -181 89 -135 136
rect -181 55 -175 89
rect -141 55 -135 89
rect -181 17 -135 55
rect -181 -17 -175 17
rect -141 -17 -135 17
rect -181 -64 -135 -17
rect -23 89 23 136
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -64 23 -17
rect 135 89 181 136
rect 135 55 141 89
rect 175 55 181 89
rect 135 17 181 55
rect 135 -17 141 17
rect 175 -17 181 17
rect 135 -64 181 -17
rect -125 -111 -33 -105
rect -125 -145 -96 -111
rect -62 -145 -33 -111
rect -125 -151 -33 -145
rect 33 -111 125 -105
rect 33 -145 62 -111
rect 96 -145 125 -111
rect 33 -151 125 -145
<< properties >>
string FIXED_BBOX -292 -267 292 267
<< end >>
