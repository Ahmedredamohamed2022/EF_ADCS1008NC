magic
tech sky130A
magscale 1 2
timestamp 1694031861
<< dnwell >>
rect -4467 -3821 2737 6561
<< nwell >>
rect -4547 6326 2817 6641
rect -4547 -3586 -4232 6326
rect 2502 -3586 2817 6326
rect -4547 -3901 2817 -3586
<< mvnsubdiff >>
rect -4481 6555 2751 6575
rect -4481 6521 -4384 6555
rect -4350 6521 -4316 6555
rect -4282 6521 -4248 6555
rect -4214 6521 -4180 6555
rect -4146 6521 -4112 6555
rect -4078 6521 -4044 6555
rect -4010 6521 -3976 6555
rect -3942 6521 -3908 6555
rect -3874 6521 -3840 6555
rect -3806 6521 -3772 6555
rect -3738 6521 -3704 6555
rect -3670 6521 -3636 6555
rect -3602 6521 -3568 6555
rect -3534 6521 -3500 6555
rect -3466 6521 -3432 6555
rect -3398 6521 -3364 6555
rect -3330 6521 -3296 6555
rect -3262 6521 -3228 6555
rect -3194 6521 -3160 6555
rect -3126 6521 -3092 6555
rect -3058 6521 -3024 6555
rect -2990 6521 -2956 6555
rect -2922 6521 -2888 6555
rect -2854 6521 -2820 6555
rect -2786 6521 -2752 6555
rect -2718 6521 -2684 6555
rect -2650 6521 -2616 6555
rect -2582 6521 -2548 6555
rect -2514 6521 -2480 6555
rect -2446 6521 -2412 6555
rect -2378 6521 -2344 6555
rect -2310 6521 -2276 6555
rect -2242 6521 -2208 6555
rect -2174 6521 -2140 6555
rect -2106 6521 -2072 6555
rect -2038 6521 -2004 6555
rect -1970 6521 -1936 6555
rect -1902 6521 -1868 6555
rect -1834 6521 -1800 6555
rect -1766 6521 -1732 6555
rect -1698 6521 -1664 6555
rect -1630 6521 -1596 6555
rect -1562 6521 -1528 6555
rect -1494 6521 -1460 6555
rect -1426 6521 -1392 6555
rect -1358 6521 -1324 6555
rect -1290 6521 -1256 6555
rect -1222 6521 -1188 6555
rect -1154 6521 -1120 6555
rect -1086 6521 -1052 6555
rect -1018 6521 -984 6555
rect -950 6521 -916 6555
rect -882 6521 -848 6555
rect -814 6521 -780 6555
rect -746 6521 -712 6555
rect -678 6521 -644 6555
rect -610 6521 -576 6555
rect -542 6521 -508 6555
rect -474 6521 -440 6555
rect -406 6521 -372 6555
rect -338 6521 -304 6555
rect -270 6521 -236 6555
rect -202 6521 -168 6555
rect -134 6521 -100 6555
rect -66 6521 -32 6555
rect 2 6521 36 6555
rect 70 6521 104 6555
rect 138 6521 172 6555
rect 206 6521 240 6555
rect 274 6521 308 6555
rect 342 6521 376 6555
rect 410 6521 444 6555
rect 478 6521 512 6555
rect 546 6521 580 6555
rect 614 6521 648 6555
rect 682 6521 716 6555
rect 750 6521 784 6555
rect 818 6521 852 6555
rect 886 6521 920 6555
rect 954 6521 988 6555
rect 1022 6521 1056 6555
rect 1090 6521 1124 6555
rect 1158 6521 1192 6555
rect 1226 6521 1260 6555
rect 1294 6521 1328 6555
rect 1362 6521 1396 6555
rect 1430 6521 1464 6555
rect 1498 6521 1532 6555
rect 1566 6521 1600 6555
rect 1634 6521 1668 6555
rect 1702 6521 1736 6555
rect 1770 6521 1804 6555
rect 1838 6521 1872 6555
rect 1906 6521 1940 6555
rect 1974 6521 2008 6555
rect 2042 6521 2076 6555
rect 2110 6521 2144 6555
rect 2178 6521 2212 6555
rect 2246 6521 2280 6555
rect 2314 6521 2348 6555
rect 2382 6521 2416 6555
rect 2450 6521 2484 6555
rect 2518 6521 2552 6555
rect 2586 6521 2620 6555
rect 2654 6521 2751 6555
rect -4481 6501 2751 6521
rect -4481 6487 -4407 6501
rect -4481 6453 -4461 6487
rect -4427 6453 -4407 6487
rect -4481 6419 -4407 6453
rect -4481 6385 -4461 6419
rect -4427 6385 -4407 6419
rect -4481 6351 -4407 6385
rect -4481 6317 -4461 6351
rect -4427 6317 -4407 6351
rect -4481 6283 -4407 6317
rect -4481 6249 -4461 6283
rect -4427 6249 -4407 6283
rect -4481 6215 -4407 6249
rect -4481 6181 -4461 6215
rect -4427 6181 -4407 6215
rect -4481 6147 -4407 6181
rect -4481 6113 -4461 6147
rect -4427 6113 -4407 6147
rect -4481 6079 -4407 6113
rect -4481 6045 -4461 6079
rect -4427 6045 -4407 6079
rect -4481 6011 -4407 6045
rect -4481 5977 -4461 6011
rect -4427 5977 -4407 6011
rect -4481 5943 -4407 5977
rect -4481 5909 -4461 5943
rect -4427 5909 -4407 5943
rect -4481 5875 -4407 5909
rect -4481 5841 -4461 5875
rect -4427 5841 -4407 5875
rect -4481 5807 -4407 5841
rect -4481 5773 -4461 5807
rect -4427 5773 -4407 5807
rect -4481 5739 -4407 5773
rect -4481 5705 -4461 5739
rect -4427 5705 -4407 5739
rect -4481 5671 -4407 5705
rect -4481 5637 -4461 5671
rect -4427 5637 -4407 5671
rect -4481 5603 -4407 5637
rect -4481 5569 -4461 5603
rect -4427 5569 -4407 5603
rect -4481 5535 -4407 5569
rect -4481 5501 -4461 5535
rect -4427 5501 -4407 5535
rect -4481 5467 -4407 5501
rect -4481 5433 -4461 5467
rect -4427 5433 -4407 5467
rect -4481 5399 -4407 5433
rect -4481 5365 -4461 5399
rect -4427 5365 -4407 5399
rect -4481 5331 -4407 5365
rect -4481 5297 -4461 5331
rect -4427 5297 -4407 5331
rect -4481 5263 -4407 5297
rect -4481 5229 -4461 5263
rect -4427 5229 -4407 5263
rect -4481 5195 -4407 5229
rect -4481 5161 -4461 5195
rect -4427 5161 -4407 5195
rect -4481 5127 -4407 5161
rect -4481 5093 -4461 5127
rect -4427 5093 -4407 5127
rect -4481 5059 -4407 5093
rect -4481 5025 -4461 5059
rect -4427 5025 -4407 5059
rect -4481 4991 -4407 5025
rect -4481 4957 -4461 4991
rect -4427 4957 -4407 4991
rect -4481 4923 -4407 4957
rect -4481 4889 -4461 4923
rect -4427 4889 -4407 4923
rect -4481 4855 -4407 4889
rect -4481 4821 -4461 4855
rect -4427 4821 -4407 4855
rect -4481 4787 -4407 4821
rect -4481 4753 -4461 4787
rect -4427 4753 -4407 4787
rect -4481 4719 -4407 4753
rect -4481 4685 -4461 4719
rect -4427 4685 -4407 4719
rect -4481 4651 -4407 4685
rect -4481 4617 -4461 4651
rect -4427 4617 -4407 4651
rect -4481 4583 -4407 4617
rect -4481 4549 -4461 4583
rect -4427 4549 -4407 4583
rect -4481 4515 -4407 4549
rect -4481 4481 -4461 4515
rect -4427 4481 -4407 4515
rect -4481 4447 -4407 4481
rect -4481 4413 -4461 4447
rect -4427 4413 -4407 4447
rect -4481 4379 -4407 4413
rect -4481 4345 -4461 4379
rect -4427 4345 -4407 4379
rect -4481 4311 -4407 4345
rect -4481 4277 -4461 4311
rect -4427 4277 -4407 4311
rect -4481 4243 -4407 4277
rect -4481 4209 -4461 4243
rect -4427 4209 -4407 4243
rect -4481 4175 -4407 4209
rect -4481 4141 -4461 4175
rect -4427 4141 -4407 4175
rect -4481 4107 -4407 4141
rect -4481 4073 -4461 4107
rect -4427 4073 -4407 4107
rect -4481 4039 -4407 4073
rect -4481 4005 -4461 4039
rect -4427 4005 -4407 4039
rect -4481 3971 -4407 4005
rect -4481 3937 -4461 3971
rect -4427 3937 -4407 3971
rect -4481 3903 -4407 3937
rect -4481 3869 -4461 3903
rect -4427 3869 -4407 3903
rect -4481 3835 -4407 3869
rect -4481 3801 -4461 3835
rect -4427 3801 -4407 3835
rect -4481 3767 -4407 3801
rect -4481 3733 -4461 3767
rect -4427 3733 -4407 3767
rect -4481 3699 -4407 3733
rect -4481 3665 -4461 3699
rect -4427 3665 -4407 3699
rect -4481 3631 -4407 3665
rect -4481 3597 -4461 3631
rect -4427 3597 -4407 3631
rect -4481 3563 -4407 3597
rect -4481 3529 -4461 3563
rect -4427 3529 -4407 3563
rect -4481 3495 -4407 3529
rect -4481 3461 -4461 3495
rect -4427 3461 -4407 3495
rect -4481 3427 -4407 3461
rect -4481 3393 -4461 3427
rect -4427 3393 -4407 3427
rect -4481 3359 -4407 3393
rect -4481 3325 -4461 3359
rect -4427 3325 -4407 3359
rect -4481 3291 -4407 3325
rect -4481 3257 -4461 3291
rect -4427 3257 -4407 3291
rect -4481 3223 -4407 3257
rect -4481 3189 -4461 3223
rect -4427 3189 -4407 3223
rect -4481 3155 -4407 3189
rect -4481 3121 -4461 3155
rect -4427 3121 -4407 3155
rect -4481 3087 -4407 3121
rect -4481 3053 -4461 3087
rect -4427 3053 -4407 3087
rect -4481 3019 -4407 3053
rect -4481 2985 -4461 3019
rect -4427 2985 -4407 3019
rect -4481 2951 -4407 2985
rect -4481 2917 -4461 2951
rect -4427 2917 -4407 2951
rect -4481 2883 -4407 2917
rect -4481 2849 -4461 2883
rect -4427 2849 -4407 2883
rect -4481 2815 -4407 2849
rect -4481 2781 -4461 2815
rect -4427 2781 -4407 2815
rect -4481 2747 -4407 2781
rect -4481 2713 -4461 2747
rect -4427 2713 -4407 2747
rect -4481 2679 -4407 2713
rect -4481 2645 -4461 2679
rect -4427 2645 -4407 2679
rect -4481 2611 -4407 2645
rect -4481 2577 -4461 2611
rect -4427 2577 -4407 2611
rect -4481 2543 -4407 2577
rect -4481 2509 -4461 2543
rect -4427 2509 -4407 2543
rect -4481 2475 -4407 2509
rect -4481 2441 -4461 2475
rect -4427 2441 -4407 2475
rect -4481 2407 -4407 2441
rect -4481 2373 -4461 2407
rect -4427 2373 -4407 2407
rect -4481 2339 -4407 2373
rect -4481 2305 -4461 2339
rect -4427 2305 -4407 2339
rect -4481 2271 -4407 2305
rect -4481 2237 -4461 2271
rect -4427 2237 -4407 2271
rect -4481 2203 -4407 2237
rect -4481 2169 -4461 2203
rect -4427 2169 -4407 2203
rect -4481 2135 -4407 2169
rect -4481 2101 -4461 2135
rect -4427 2101 -4407 2135
rect -4481 2067 -4407 2101
rect -4481 2033 -4461 2067
rect -4427 2033 -4407 2067
rect -4481 1999 -4407 2033
rect -4481 1965 -4461 1999
rect -4427 1965 -4407 1999
rect -4481 1931 -4407 1965
rect -4481 1897 -4461 1931
rect -4427 1897 -4407 1931
rect -4481 1863 -4407 1897
rect -4481 1829 -4461 1863
rect -4427 1829 -4407 1863
rect -4481 1795 -4407 1829
rect -4481 1761 -4461 1795
rect -4427 1761 -4407 1795
rect -4481 1727 -4407 1761
rect -4481 1693 -4461 1727
rect -4427 1693 -4407 1727
rect -4481 1659 -4407 1693
rect -4481 1625 -4461 1659
rect -4427 1625 -4407 1659
rect -4481 1591 -4407 1625
rect -4481 1557 -4461 1591
rect -4427 1557 -4407 1591
rect -4481 1523 -4407 1557
rect -4481 1489 -4461 1523
rect -4427 1489 -4407 1523
rect -4481 1455 -4407 1489
rect -4481 1421 -4461 1455
rect -4427 1421 -4407 1455
rect -4481 1387 -4407 1421
rect -4481 1353 -4461 1387
rect -4427 1353 -4407 1387
rect -4481 1319 -4407 1353
rect -4481 1285 -4461 1319
rect -4427 1285 -4407 1319
rect -4481 1251 -4407 1285
rect -4481 1217 -4461 1251
rect -4427 1217 -4407 1251
rect -4481 1183 -4407 1217
rect -4481 1149 -4461 1183
rect -4427 1149 -4407 1183
rect -4481 1115 -4407 1149
rect -4481 1081 -4461 1115
rect -4427 1081 -4407 1115
rect -4481 1047 -4407 1081
rect -4481 1013 -4461 1047
rect -4427 1013 -4407 1047
rect -4481 979 -4407 1013
rect -4481 945 -4461 979
rect -4427 945 -4407 979
rect -4481 911 -4407 945
rect -4481 877 -4461 911
rect -4427 877 -4407 911
rect -4481 843 -4407 877
rect -4481 809 -4461 843
rect -4427 809 -4407 843
rect -4481 775 -4407 809
rect -4481 741 -4461 775
rect -4427 741 -4407 775
rect -4481 707 -4407 741
rect -4481 673 -4461 707
rect -4427 673 -4407 707
rect -4481 639 -4407 673
rect -4481 605 -4461 639
rect -4427 605 -4407 639
rect -4481 571 -4407 605
rect -4481 537 -4461 571
rect -4427 537 -4407 571
rect -4481 503 -4407 537
rect -4481 469 -4461 503
rect -4427 469 -4407 503
rect -4481 435 -4407 469
rect -4481 401 -4461 435
rect -4427 401 -4407 435
rect -4481 367 -4407 401
rect -4481 333 -4461 367
rect -4427 333 -4407 367
rect -4481 299 -4407 333
rect -4481 265 -4461 299
rect -4427 265 -4407 299
rect -4481 231 -4407 265
rect -4481 197 -4461 231
rect -4427 197 -4407 231
rect -4481 163 -4407 197
rect -4481 129 -4461 163
rect -4427 129 -4407 163
rect -4481 95 -4407 129
rect -4481 61 -4461 95
rect -4427 61 -4407 95
rect -4481 27 -4407 61
rect -4481 -7 -4461 27
rect -4427 -7 -4407 27
rect -4481 -41 -4407 -7
rect -4481 -75 -4461 -41
rect -4427 -75 -4407 -41
rect -4481 -109 -4407 -75
rect -4481 -143 -4461 -109
rect -4427 -143 -4407 -109
rect -4481 -177 -4407 -143
rect -4481 -211 -4461 -177
rect -4427 -211 -4407 -177
rect -4481 -245 -4407 -211
rect -4481 -279 -4461 -245
rect -4427 -279 -4407 -245
rect -4481 -313 -4407 -279
rect -4481 -347 -4461 -313
rect -4427 -347 -4407 -313
rect -4481 -381 -4407 -347
rect -4481 -415 -4461 -381
rect -4427 -415 -4407 -381
rect -4481 -449 -4407 -415
rect -4481 -483 -4461 -449
rect -4427 -483 -4407 -449
rect -4481 -517 -4407 -483
rect -4481 -551 -4461 -517
rect -4427 -551 -4407 -517
rect -4481 -585 -4407 -551
rect -4481 -619 -4461 -585
rect -4427 -619 -4407 -585
rect -4481 -653 -4407 -619
rect -4481 -687 -4461 -653
rect -4427 -687 -4407 -653
rect -4481 -721 -4407 -687
rect -4481 -755 -4461 -721
rect -4427 -755 -4407 -721
rect -4481 -789 -4407 -755
rect -4481 -823 -4461 -789
rect -4427 -823 -4407 -789
rect -4481 -857 -4407 -823
rect -4481 -891 -4461 -857
rect -4427 -891 -4407 -857
rect -4481 -925 -4407 -891
rect -4481 -959 -4461 -925
rect -4427 -959 -4407 -925
rect -4481 -993 -4407 -959
rect -4481 -1027 -4461 -993
rect -4427 -1027 -4407 -993
rect -4481 -1061 -4407 -1027
rect -4481 -1095 -4461 -1061
rect -4427 -1095 -4407 -1061
rect -4481 -1129 -4407 -1095
rect -4481 -1163 -4461 -1129
rect -4427 -1163 -4407 -1129
rect -4481 -1197 -4407 -1163
rect -4481 -1231 -4461 -1197
rect -4427 -1231 -4407 -1197
rect -4481 -1265 -4407 -1231
rect -4481 -1299 -4461 -1265
rect -4427 -1299 -4407 -1265
rect -4481 -1333 -4407 -1299
rect -4481 -1367 -4461 -1333
rect -4427 -1367 -4407 -1333
rect -4481 -1401 -4407 -1367
rect -4481 -1435 -4461 -1401
rect -4427 -1435 -4407 -1401
rect -4481 -1469 -4407 -1435
rect -4481 -1503 -4461 -1469
rect -4427 -1503 -4407 -1469
rect -4481 -1537 -4407 -1503
rect -4481 -1571 -4461 -1537
rect -4427 -1571 -4407 -1537
rect -4481 -1605 -4407 -1571
rect -4481 -1639 -4461 -1605
rect -4427 -1639 -4407 -1605
rect -4481 -1673 -4407 -1639
rect -4481 -1707 -4461 -1673
rect -4427 -1707 -4407 -1673
rect -4481 -1741 -4407 -1707
rect -4481 -1775 -4461 -1741
rect -4427 -1775 -4407 -1741
rect -4481 -1809 -4407 -1775
rect -4481 -1843 -4461 -1809
rect -4427 -1843 -4407 -1809
rect -4481 -1877 -4407 -1843
rect -4481 -1911 -4461 -1877
rect -4427 -1911 -4407 -1877
rect -4481 -1945 -4407 -1911
rect -4481 -1979 -4461 -1945
rect -4427 -1979 -4407 -1945
rect -4481 -2013 -4407 -1979
rect -4481 -2047 -4461 -2013
rect -4427 -2047 -4407 -2013
rect -4481 -2081 -4407 -2047
rect -4481 -2115 -4461 -2081
rect -4427 -2115 -4407 -2081
rect -4481 -2149 -4407 -2115
rect -4481 -2183 -4461 -2149
rect -4427 -2183 -4407 -2149
rect -4481 -2217 -4407 -2183
rect -4481 -2251 -4461 -2217
rect -4427 -2251 -4407 -2217
rect -4481 -2285 -4407 -2251
rect -4481 -2319 -4461 -2285
rect -4427 -2319 -4407 -2285
rect -4481 -2353 -4407 -2319
rect -4481 -2387 -4461 -2353
rect -4427 -2387 -4407 -2353
rect -4481 -2421 -4407 -2387
rect -4481 -2455 -4461 -2421
rect -4427 -2455 -4407 -2421
rect -4481 -2489 -4407 -2455
rect -4481 -2523 -4461 -2489
rect -4427 -2523 -4407 -2489
rect -4481 -2557 -4407 -2523
rect -4481 -2591 -4461 -2557
rect -4427 -2591 -4407 -2557
rect -4481 -2625 -4407 -2591
rect -4481 -2659 -4461 -2625
rect -4427 -2659 -4407 -2625
rect -4481 -2693 -4407 -2659
rect -4481 -2727 -4461 -2693
rect -4427 -2727 -4407 -2693
rect -4481 -2761 -4407 -2727
rect -4481 -2795 -4461 -2761
rect -4427 -2795 -4407 -2761
rect -4481 -2829 -4407 -2795
rect -4481 -2863 -4461 -2829
rect -4427 -2863 -4407 -2829
rect -4481 -2897 -4407 -2863
rect -4481 -2931 -4461 -2897
rect -4427 -2931 -4407 -2897
rect -4481 -2965 -4407 -2931
rect -4481 -2999 -4461 -2965
rect -4427 -2999 -4407 -2965
rect -4481 -3033 -4407 -2999
rect -4481 -3067 -4461 -3033
rect -4427 -3067 -4407 -3033
rect -4481 -3101 -4407 -3067
rect -4481 -3135 -4461 -3101
rect -4427 -3135 -4407 -3101
rect -4481 -3169 -4407 -3135
rect -4481 -3203 -4461 -3169
rect -4427 -3203 -4407 -3169
rect -4481 -3237 -4407 -3203
rect -4481 -3271 -4461 -3237
rect -4427 -3271 -4407 -3237
rect -4481 -3305 -4407 -3271
rect -4481 -3339 -4461 -3305
rect -4427 -3339 -4407 -3305
rect -4481 -3373 -4407 -3339
rect -4481 -3407 -4461 -3373
rect -4427 -3407 -4407 -3373
rect -4481 -3441 -4407 -3407
rect -4481 -3475 -4461 -3441
rect -4427 -3475 -4407 -3441
rect -4481 -3509 -4407 -3475
rect -4481 -3543 -4461 -3509
rect -4427 -3543 -4407 -3509
rect -4481 -3577 -4407 -3543
rect -4481 -3611 -4461 -3577
rect -4427 -3611 -4407 -3577
rect -4481 -3645 -4407 -3611
rect -4481 -3679 -4461 -3645
rect -4427 -3679 -4407 -3645
rect -4481 -3713 -4407 -3679
rect -4481 -3747 -4461 -3713
rect -4427 -3747 -4407 -3713
rect -4481 -3761 -4407 -3747
rect 2677 6487 2751 6501
rect 2677 6453 2697 6487
rect 2731 6453 2751 6487
rect 2677 6419 2751 6453
rect 2677 6385 2697 6419
rect 2731 6385 2751 6419
rect 2677 6351 2751 6385
rect 2677 6317 2697 6351
rect 2731 6317 2751 6351
rect 2677 6283 2751 6317
rect 2677 6249 2697 6283
rect 2731 6249 2751 6283
rect 2677 6215 2751 6249
rect 2677 6181 2697 6215
rect 2731 6181 2751 6215
rect 2677 6147 2751 6181
rect 2677 6113 2697 6147
rect 2731 6113 2751 6147
rect 2677 6079 2751 6113
rect 2677 6045 2697 6079
rect 2731 6045 2751 6079
rect 2677 6011 2751 6045
rect 2677 5977 2697 6011
rect 2731 5977 2751 6011
rect 2677 5943 2751 5977
rect 2677 5909 2697 5943
rect 2731 5909 2751 5943
rect 2677 5875 2751 5909
rect 2677 5841 2697 5875
rect 2731 5841 2751 5875
rect 2677 5807 2751 5841
rect 2677 5773 2697 5807
rect 2731 5773 2751 5807
rect 2677 5739 2751 5773
rect 2677 5705 2697 5739
rect 2731 5705 2751 5739
rect 2677 5671 2751 5705
rect 2677 5637 2697 5671
rect 2731 5637 2751 5671
rect 2677 5603 2751 5637
rect 2677 5569 2697 5603
rect 2731 5569 2751 5603
rect 2677 5535 2751 5569
rect 2677 5501 2697 5535
rect 2731 5501 2751 5535
rect 2677 5467 2751 5501
rect 2677 5433 2697 5467
rect 2731 5433 2751 5467
rect 2677 5399 2751 5433
rect 2677 5365 2697 5399
rect 2731 5365 2751 5399
rect 2677 5331 2751 5365
rect 2677 5297 2697 5331
rect 2731 5297 2751 5331
rect 2677 5263 2751 5297
rect 2677 5229 2697 5263
rect 2731 5229 2751 5263
rect 2677 5195 2751 5229
rect 2677 5161 2697 5195
rect 2731 5161 2751 5195
rect 2677 5127 2751 5161
rect 2677 5093 2697 5127
rect 2731 5093 2751 5127
rect 2677 5059 2751 5093
rect 2677 5025 2697 5059
rect 2731 5025 2751 5059
rect 2677 4991 2751 5025
rect 2677 4957 2697 4991
rect 2731 4957 2751 4991
rect 2677 4923 2751 4957
rect 2677 4889 2697 4923
rect 2731 4889 2751 4923
rect 2677 4855 2751 4889
rect 2677 4821 2697 4855
rect 2731 4821 2751 4855
rect 2677 4787 2751 4821
rect 2677 4753 2697 4787
rect 2731 4753 2751 4787
rect 2677 4719 2751 4753
rect 2677 4685 2697 4719
rect 2731 4685 2751 4719
rect 2677 4651 2751 4685
rect 2677 4617 2697 4651
rect 2731 4617 2751 4651
rect 2677 4583 2751 4617
rect 2677 4549 2697 4583
rect 2731 4549 2751 4583
rect 2677 4515 2751 4549
rect 2677 4481 2697 4515
rect 2731 4481 2751 4515
rect 2677 4447 2751 4481
rect 2677 4413 2697 4447
rect 2731 4413 2751 4447
rect 2677 4379 2751 4413
rect 2677 4345 2697 4379
rect 2731 4345 2751 4379
rect 2677 4311 2751 4345
rect 2677 4277 2697 4311
rect 2731 4277 2751 4311
rect 2677 4243 2751 4277
rect 2677 4209 2697 4243
rect 2731 4209 2751 4243
rect 2677 4175 2751 4209
rect 2677 4141 2697 4175
rect 2731 4141 2751 4175
rect 2677 4107 2751 4141
rect 2677 4073 2697 4107
rect 2731 4073 2751 4107
rect 2677 4039 2751 4073
rect 2677 4005 2697 4039
rect 2731 4005 2751 4039
rect 2677 3971 2751 4005
rect 2677 3937 2697 3971
rect 2731 3937 2751 3971
rect 2677 3903 2751 3937
rect 2677 3869 2697 3903
rect 2731 3869 2751 3903
rect 2677 3835 2751 3869
rect 2677 3801 2697 3835
rect 2731 3801 2751 3835
rect 2677 3767 2751 3801
rect 2677 3733 2697 3767
rect 2731 3733 2751 3767
rect 2677 3699 2751 3733
rect 2677 3665 2697 3699
rect 2731 3665 2751 3699
rect 2677 3631 2751 3665
rect 2677 3597 2697 3631
rect 2731 3597 2751 3631
rect 2677 3563 2751 3597
rect 2677 3529 2697 3563
rect 2731 3529 2751 3563
rect 2677 3495 2751 3529
rect 2677 3461 2697 3495
rect 2731 3461 2751 3495
rect 2677 3427 2751 3461
rect 2677 3393 2697 3427
rect 2731 3393 2751 3427
rect 2677 3359 2751 3393
rect 2677 3325 2697 3359
rect 2731 3325 2751 3359
rect 2677 3291 2751 3325
rect 2677 3257 2697 3291
rect 2731 3257 2751 3291
rect 2677 3223 2751 3257
rect 2677 3189 2697 3223
rect 2731 3189 2751 3223
rect 2677 3155 2751 3189
rect 2677 3121 2697 3155
rect 2731 3121 2751 3155
rect 2677 3087 2751 3121
rect 2677 3053 2697 3087
rect 2731 3053 2751 3087
rect 2677 3019 2751 3053
rect 2677 2985 2697 3019
rect 2731 2985 2751 3019
rect 2677 2951 2751 2985
rect 2677 2917 2697 2951
rect 2731 2917 2751 2951
rect 2677 2883 2751 2917
rect 2677 2849 2697 2883
rect 2731 2849 2751 2883
rect 2677 2815 2751 2849
rect 2677 2781 2697 2815
rect 2731 2781 2751 2815
rect 2677 2747 2751 2781
rect 2677 2713 2697 2747
rect 2731 2713 2751 2747
rect 2677 2679 2751 2713
rect 2677 2645 2697 2679
rect 2731 2645 2751 2679
rect 2677 2611 2751 2645
rect 2677 2577 2697 2611
rect 2731 2577 2751 2611
rect 2677 2543 2751 2577
rect 2677 2509 2697 2543
rect 2731 2509 2751 2543
rect 2677 2475 2751 2509
rect 2677 2441 2697 2475
rect 2731 2441 2751 2475
rect 2677 2407 2751 2441
rect 2677 2373 2697 2407
rect 2731 2373 2751 2407
rect 2677 2339 2751 2373
rect 2677 2305 2697 2339
rect 2731 2305 2751 2339
rect 2677 2271 2751 2305
rect 2677 2237 2697 2271
rect 2731 2237 2751 2271
rect 2677 2203 2751 2237
rect 2677 2169 2697 2203
rect 2731 2169 2751 2203
rect 2677 2135 2751 2169
rect 2677 2101 2697 2135
rect 2731 2101 2751 2135
rect 2677 2067 2751 2101
rect 2677 2033 2697 2067
rect 2731 2033 2751 2067
rect 2677 1999 2751 2033
rect 2677 1965 2697 1999
rect 2731 1965 2751 1999
rect 2677 1931 2751 1965
rect 2677 1897 2697 1931
rect 2731 1897 2751 1931
rect 2677 1863 2751 1897
rect 2677 1829 2697 1863
rect 2731 1829 2751 1863
rect 2677 1795 2751 1829
rect 2677 1761 2697 1795
rect 2731 1761 2751 1795
rect 2677 1727 2751 1761
rect 2677 1693 2697 1727
rect 2731 1693 2751 1727
rect 2677 1659 2751 1693
rect 2677 1625 2697 1659
rect 2731 1625 2751 1659
rect 2677 1591 2751 1625
rect 2677 1557 2697 1591
rect 2731 1557 2751 1591
rect 2677 1523 2751 1557
rect 2677 1489 2697 1523
rect 2731 1489 2751 1523
rect 2677 1455 2751 1489
rect 2677 1421 2697 1455
rect 2731 1421 2751 1455
rect 2677 1387 2751 1421
rect 2677 1353 2697 1387
rect 2731 1353 2751 1387
rect 2677 1319 2751 1353
rect 2677 1285 2697 1319
rect 2731 1285 2751 1319
rect 2677 1251 2751 1285
rect 2677 1217 2697 1251
rect 2731 1217 2751 1251
rect 2677 1183 2751 1217
rect 2677 1149 2697 1183
rect 2731 1149 2751 1183
rect 2677 1115 2751 1149
rect 2677 1081 2697 1115
rect 2731 1081 2751 1115
rect 2677 1047 2751 1081
rect 2677 1013 2697 1047
rect 2731 1013 2751 1047
rect 2677 979 2751 1013
rect 2677 945 2697 979
rect 2731 945 2751 979
rect 2677 911 2751 945
rect 2677 877 2697 911
rect 2731 877 2751 911
rect 2677 843 2751 877
rect 2677 809 2697 843
rect 2731 809 2751 843
rect 2677 775 2751 809
rect 2677 741 2697 775
rect 2731 741 2751 775
rect 2677 707 2751 741
rect 2677 673 2697 707
rect 2731 673 2751 707
rect 2677 639 2751 673
rect 2677 605 2697 639
rect 2731 605 2751 639
rect 2677 571 2751 605
rect 2677 537 2697 571
rect 2731 537 2751 571
rect 2677 503 2751 537
rect 2677 469 2697 503
rect 2731 469 2751 503
rect 2677 435 2751 469
rect 2677 401 2697 435
rect 2731 401 2751 435
rect 2677 367 2751 401
rect 2677 333 2697 367
rect 2731 333 2751 367
rect 2677 299 2751 333
rect 2677 265 2697 299
rect 2731 265 2751 299
rect 2677 231 2751 265
rect 2677 197 2697 231
rect 2731 197 2751 231
rect 2677 163 2751 197
rect 2677 129 2697 163
rect 2731 129 2751 163
rect 2677 95 2751 129
rect 2677 61 2697 95
rect 2731 61 2751 95
rect 2677 27 2751 61
rect 2677 -7 2697 27
rect 2731 -7 2751 27
rect 2677 -41 2751 -7
rect 2677 -75 2697 -41
rect 2731 -75 2751 -41
rect 2677 -109 2751 -75
rect 2677 -143 2697 -109
rect 2731 -143 2751 -109
rect 2677 -177 2751 -143
rect 2677 -211 2697 -177
rect 2731 -211 2751 -177
rect 2677 -245 2751 -211
rect 2677 -279 2697 -245
rect 2731 -279 2751 -245
rect 2677 -313 2751 -279
rect 2677 -347 2697 -313
rect 2731 -347 2751 -313
rect 2677 -381 2751 -347
rect 2677 -415 2697 -381
rect 2731 -415 2751 -381
rect 2677 -449 2751 -415
rect 2677 -483 2697 -449
rect 2731 -483 2751 -449
rect 2677 -517 2751 -483
rect 2677 -551 2697 -517
rect 2731 -551 2751 -517
rect 2677 -585 2751 -551
rect 2677 -619 2697 -585
rect 2731 -619 2751 -585
rect 2677 -653 2751 -619
rect 2677 -687 2697 -653
rect 2731 -687 2751 -653
rect 2677 -721 2751 -687
rect 2677 -755 2697 -721
rect 2731 -755 2751 -721
rect 2677 -789 2751 -755
rect 2677 -823 2697 -789
rect 2731 -823 2751 -789
rect 2677 -857 2751 -823
rect 2677 -891 2697 -857
rect 2731 -891 2751 -857
rect 2677 -925 2751 -891
rect 2677 -959 2697 -925
rect 2731 -959 2751 -925
rect 2677 -993 2751 -959
rect 2677 -1027 2697 -993
rect 2731 -1027 2751 -993
rect 2677 -1061 2751 -1027
rect 2677 -1095 2697 -1061
rect 2731 -1095 2751 -1061
rect 2677 -1129 2751 -1095
rect 2677 -1163 2697 -1129
rect 2731 -1163 2751 -1129
rect 2677 -1197 2751 -1163
rect 2677 -1231 2697 -1197
rect 2731 -1231 2751 -1197
rect 2677 -1265 2751 -1231
rect 2677 -1299 2697 -1265
rect 2731 -1299 2751 -1265
rect 2677 -1333 2751 -1299
rect 2677 -1367 2697 -1333
rect 2731 -1367 2751 -1333
rect 2677 -1401 2751 -1367
rect 2677 -1435 2697 -1401
rect 2731 -1435 2751 -1401
rect 2677 -1469 2751 -1435
rect 2677 -1503 2697 -1469
rect 2731 -1503 2751 -1469
rect 2677 -1537 2751 -1503
rect 2677 -1571 2697 -1537
rect 2731 -1571 2751 -1537
rect 2677 -1605 2751 -1571
rect 2677 -1639 2697 -1605
rect 2731 -1639 2751 -1605
rect 2677 -1673 2751 -1639
rect 2677 -1707 2697 -1673
rect 2731 -1707 2751 -1673
rect 2677 -1741 2751 -1707
rect 2677 -1775 2697 -1741
rect 2731 -1775 2751 -1741
rect 2677 -1809 2751 -1775
rect 2677 -1843 2697 -1809
rect 2731 -1843 2751 -1809
rect 2677 -1877 2751 -1843
rect 2677 -1911 2697 -1877
rect 2731 -1911 2751 -1877
rect 2677 -1945 2751 -1911
rect 2677 -1979 2697 -1945
rect 2731 -1979 2751 -1945
rect 2677 -2013 2751 -1979
rect 2677 -2047 2697 -2013
rect 2731 -2047 2751 -2013
rect 2677 -2081 2751 -2047
rect 2677 -2115 2697 -2081
rect 2731 -2115 2751 -2081
rect 2677 -2149 2751 -2115
rect 2677 -2183 2697 -2149
rect 2731 -2183 2751 -2149
rect 2677 -2217 2751 -2183
rect 2677 -2251 2697 -2217
rect 2731 -2251 2751 -2217
rect 2677 -2285 2751 -2251
rect 2677 -2319 2697 -2285
rect 2731 -2319 2751 -2285
rect 2677 -2353 2751 -2319
rect 2677 -2387 2697 -2353
rect 2731 -2387 2751 -2353
rect 2677 -2421 2751 -2387
rect 2677 -2455 2697 -2421
rect 2731 -2455 2751 -2421
rect 2677 -2489 2751 -2455
rect 2677 -2523 2697 -2489
rect 2731 -2523 2751 -2489
rect 2677 -2557 2751 -2523
rect 2677 -2591 2697 -2557
rect 2731 -2591 2751 -2557
rect 2677 -2625 2751 -2591
rect 2677 -2659 2697 -2625
rect 2731 -2659 2751 -2625
rect 2677 -2693 2751 -2659
rect 2677 -2727 2697 -2693
rect 2731 -2727 2751 -2693
rect 2677 -2761 2751 -2727
rect 2677 -2795 2697 -2761
rect 2731 -2795 2751 -2761
rect 2677 -2829 2751 -2795
rect 2677 -2863 2697 -2829
rect 2731 -2863 2751 -2829
rect 2677 -2897 2751 -2863
rect 2677 -2931 2697 -2897
rect 2731 -2931 2751 -2897
rect 2677 -2965 2751 -2931
rect 2677 -2999 2697 -2965
rect 2731 -2999 2751 -2965
rect 2677 -3033 2751 -2999
rect 2677 -3067 2697 -3033
rect 2731 -3067 2751 -3033
rect 2677 -3101 2751 -3067
rect 2677 -3135 2697 -3101
rect 2731 -3135 2751 -3101
rect 2677 -3169 2751 -3135
rect 2677 -3203 2697 -3169
rect 2731 -3203 2751 -3169
rect 2677 -3237 2751 -3203
rect 2677 -3271 2697 -3237
rect 2731 -3271 2751 -3237
rect 2677 -3305 2751 -3271
rect 2677 -3339 2697 -3305
rect 2731 -3339 2751 -3305
rect 2677 -3373 2751 -3339
rect 2677 -3407 2697 -3373
rect 2731 -3407 2751 -3373
rect 2677 -3441 2751 -3407
rect 2677 -3475 2697 -3441
rect 2731 -3475 2751 -3441
rect 2677 -3509 2751 -3475
rect 2677 -3543 2697 -3509
rect 2731 -3543 2751 -3509
rect 2677 -3577 2751 -3543
rect 2677 -3611 2697 -3577
rect 2731 -3611 2751 -3577
rect 2677 -3645 2751 -3611
rect 2677 -3679 2697 -3645
rect 2731 -3679 2751 -3645
rect 2677 -3713 2751 -3679
rect 2677 -3747 2697 -3713
rect 2731 -3747 2751 -3713
rect 2677 -3761 2751 -3747
rect -4481 -3781 2751 -3761
rect -4481 -3815 -4384 -3781
rect -4350 -3815 -4316 -3781
rect -4282 -3815 -4248 -3781
rect -4214 -3815 -4180 -3781
rect -4146 -3815 -4112 -3781
rect -4078 -3815 -4044 -3781
rect -4010 -3815 -3976 -3781
rect -3942 -3815 -3908 -3781
rect -3874 -3815 -3840 -3781
rect -3806 -3815 -3772 -3781
rect -3738 -3815 -3704 -3781
rect -3670 -3815 -3636 -3781
rect -3602 -3815 -3568 -3781
rect -3534 -3815 -3500 -3781
rect -3466 -3815 -3432 -3781
rect -3398 -3815 -3364 -3781
rect -3330 -3815 -3296 -3781
rect -3262 -3815 -3228 -3781
rect -3194 -3815 -3160 -3781
rect -3126 -3815 -3092 -3781
rect -3058 -3815 -3024 -3781
rect -2990 -3815 -2956 -3781
rect -2922 -3815 -2888 -3781
rect -2854 -3815 -2820 -3781
rect -2786 -3815 -2752 -3781
rect -2718 -3815 -2684 -3781
rect -2650 -3815 -2616 -3781
rect -2582 -3815 -2548 -3781
rect -2514 -3815 -2480 -3781
rect -2446 -3815 -2412 -3781
rect -2378 -3815 -2344 -3781
rect -2310 -3815 -2276 -3781
rect -2242 -3815 -2208 -3781
rect -2174 -3815 -2140 -3781
rect -2106 -3815 -2072 -3781
rect -2038 -3815 -2004 -3781
rect -1970 -3815 -1936 -3781
rect -1902 -3815 -1868 -3781
rect -1834 -3815 -1800 -3781
rect -1766 -3815 -1732 -3781
rect -1698 -3815 -1664 -3781
rect -1630 -3815 -1596 -3781
rect -1562 -3815 -1528 -3781
rect -1494 -3815 -1460 -3781
rect -1426 -3815 -1392 -3781
rect -1358 -3815 -1324 -3781
rect -1290 -3815 -1256 -3781
rect -1222 -3815 -1188 -3781
rect -1154 -3815 -1120 -3781
rect -1086 -3815 -1052 -3781
rect -1018 -3815 -984 -3781
rect -950 -3815 -916 -3781
rect -882 -3815 -848 -3781
rect -814 -3815 -780 -3781
rect -746 -3815 -712 -3781
rect -678 -3815 -644 -3781
rect -610 -3815 -576 -3781
rect -542 -3815 -508 -3781
rect -474 -3815 -440 -3781
rect -406 -3815 -372 -3781
rect -338 -3815 -304 -3781
rect -270 -3815 -236 -3781
rect -202 -3815 -168 -3781
rect -134 -3815 -100 -3781
rect -66 -3815 -32 -3781
rect 2 -3815 36 -3781
rect 70 -3815 104 -3781
rect 138 -3815 172 -3781
rect 206 -3815 240 -3781
rect 274 -3815 308 -3781
rect 342 -3815 376 -3781
rect 410 -3815 444 -3781
rect 478 -3815 512 -3781
rect 546 -3815 580 -3781
rect 614 -3815 648 -3781
rect 682 -3815 716 -3781
rect 750 -3815 784 -3781
rect 818 -3815 852 -3781
rect 886 -3815 920 -3781
rect 954 -3815 988 -3781
rect 1022 -3815 1056 -3781
rect 1090 -3815 1124 -3781
rect 1158 -3815 1192 -3781
rect 1226 -3815 1260 -3781
rect 1294 -3815 1328 -3781
rect 1362 -3815 1396 -3781
rect 1430 -3815 1464 -3781
rect 1498 -3815 1532 -3781
rect 1566 -3815 1600 -3781
rect 1634 -3815 1668 -3781
rect 1702 -3815 1736 -3781
rect 1770 -3815 1804 -3781
rect 1838 -3815 1872 -3781
rect 1906 -3815 1940 -3781
rect 1974 -3815 2008 -3781
rect 2042 -3815 2076 -3781
rect 2110 -3815 2144 -3781
rect 2178 -3815 2212 -3781
rect 2246 -3815 2280 -3781
rect 2314 -3815 2348 -3781
rect 2382 -3815 2416 -3781
rect 2450 -3815 2484 -3781
rect 2518 -3815 2552 -3781
rect 2586 -3815 2620 -3781
rect 2654 -3815 2751 -3781
rect -4481 -3835 2751 -3815
<< mvnsubdiffcont >>
rect -4384 6521 -4350 6555
rect -4316 6521 -4282 6555
rect -4248 6521 -4214 6555
rect -4180 6521 -4146 6555
rect -4112 6521 -4078 6555
rect -4044 6521 -4010 6555
rect -3976 6521 -3942 6555
rect -3908 6521 -3874 6555
rect -3840 6521 -3806 6555
rect -3772 6521 -3738 6555
rect -3704 6521 -3670 6555
rect -3636 6521 -3602 6555
rect -3568 6521 -3534 6555
rect -3500 6521 -3466 6555
rect -3432 6521 -3398 6555
rect -3364 6521 -3330 6555
rect -3296 6521 -3262 6555
rect -3228 6521 -3194 6555
rect -3160 6521 -3126 6555
rect -3092 6521 -3058 6555
rect -3024 6521 -2990 6555
rect -2956 6521 -2922 6555
rect -2888 6521 -2854 6555
rect -2820 6521 -2786 6555
rect -2752 6521 -2718 6555
rect -2684 6521 -2650 6555
rect -2616 6521 -2582 6555
rect -2548 6521 -2514 6555
rect -2480 6521 -2446 6555
rect -2412 6521 -2378 6555
rect -2344 6521 -2310 6555
rect -2276 6521 -2242 6555
rect -2208 6521 -2174 6555
rect -2140 6521 -2106 6555
rect -2072 6521 -2038 6555
rect -2004 6521 -1970 6555
rect -1936 6521 -1902 6555
rect -1868 6521 -1834 6555
rect -1800 6521 -1766 6555
rect -1732 6521 -1698 6555
rect -1664 6521 -1630 6555
rect -1596 6521 -1562 6555
rect -1528 6521 -1494 6555
rect -1460 6521 -1426 6555
rect -1392 6521 -1358 6555
rect -1324 6521 -1290 6555
rect -1256 6521 -1222 6555
rect -1188 6521 -1154 6555
rect -1120 6521 -1086 6555
rect -1052 6521 -1018 6555
rect -984 6521 -950 6555
rect -916 6521 -882 6555
rect -848 6521 -814 6555
rect -780 6521 -746 6555
rect -712 6521 -678 6555
rect -644 6521 -610 6555
rect -576 6521 -542 6555
rect -508 6521 -474 6555
rect -440 6521 -406 6555
rect -372 6521 -338 6555
rect -304 6521 -270 6555
rect -236 6521 -202 6555
rect -168 6521 -134 6555
rect -100 6521 -66 6555
rect -32 6521 2 6555
rect 36 6521 70 6555
rect 104 6521 138 6555
rect 172 6521 206 6555
rect 240 6521 274 6555
rect 308 6521 342 6555
rect 376 6521 410 6555
rect 444 6521 478 6555
rect 512 6521 546 6555
rect 580 6521 614 6555
rect 648 6521 682 6555
rect 716 6521 750 6555
rect 784 6521 818 6555
rect 852 6521 886 6555
rect 920 6521 954 6555
rect 988 6521 1022 6555
rect 1056 6521 1090 6555
rect 1124 6521 1158 6555
rect 1192 6521 1226 6555
rect 1260 6521 1294 6555
rect 1328 6521 1362 6555
rect 1396 6521 1430 6555
rect 1464 6521 1498 6555
rect 1532 6521 1566 6555
rect 1600 6521 1634 6555
rect 1668 6521 1702 6555
rect 1736 6521 1770 6555
rect 1804 6521 1838 6555
rect 1872 6521 1906 6555
rect 1940 6521 1974 6555
rect 2008 6521 2042 6555
rect 2076 6521 2110 6555
rect 2144 6521 2178 6555
rect 2212 6521 2246 6555
rect 2280 6521 2314 6555
rect 2348 6521 2382 6555
rect 2416 6521 2450 6555
rect 2484 6521 2518 6555
rect 2552 6521 2586 6555
rect 2620 6521 2654 6555
rect -4461 6453 -4427 6487
rect -4461 6385 -4427 6419
rect -4461 6317 -4427 6351
rect -4461 6249 -4427 6283
rect -4461 6181 -4427 6215
rect -4461 6113 -4427 6147
rect -4461 6045 -4427 6079
rect -4461 5977 -4427 6011
rect -4461 5909 -4427 5943
rect -4461 5841 -4427 5875
rect -4461 5773 -4427 5807
rect -4461 5705 -4427 5739
rect -4461 5637 -4427 5671
rect -4461 5569 -4427 5603
rect -4461 5501 -4427 5535
rect -4461 5433 -4427 5467
rect -4461 5365 -4427 5399
rect -4461 5297 -4427 5331
rect -4461 5229 -4427 5263
rect -4461 5161 -4427 5195
rect -4461 5093 -4427 5127
rect -4461 5025 -4427 5059
rect -4461 4957 -4427 4991
rect -4461 4889 -4427 4923
rect -4461 4821 -4427 4855
rect -4461 4753 -4427 4787
rect -4461 4685 -4427 4719
rect -4461 4617 -4427 4651
rect -4461 4549 -4427 4583
rect -4461 4481 -4427 4515
rect -4461 4413 -4427 4447
rect -4461 4345 -4427 4379
rect -4461 4277 -4427 4311
rect -4461 4209 -4427 4243
rect -4461 4141 -4427 4175
rect -4461 4073 -4427 4107
rect -4461 4005 -4427 4039
rect -4461 3937 -4427 3971
rect -4461 3869 -4427 3903
rect -4461 3801 -4427 3835
rect -4461 3733 -4427 3767
rect -4461 3665 -4427 3699
rect -4461 3597 -4427 3631
rect -4461 3529 -4427 3563
rect -4461 3461 -4427 3495
rect -4461 3393 -4427 3427
rect -4461 3325 -4427 3359
rect -4461 3257 -4427 3291
rect -4461 3189 -4427 3223
rect -4461 3121 -4427 3155
rect -4461 3053 -4427 3087
rect -4461 2985 -4427 3019
rect -4461 2917 -4427 2951
rect -4461 2849 -4427 2883
rect -4461 2781 -4427 2815
rect -4461 2713 -4427 2747
rect -4461 2645 -4427 2679
rect -4461 2577 -4427 2611
rect -4461 2509 -4427 2543
rect -4461 2441 -4427 2475
rect -4461 2373 -4427 2407
rect -4461 2305 -4427 2339
rect -4461 2237 -4427 2271
rect -4461 2169 -4427 2203
rect -4461 2101 -4427 2135
rect -4461 2033 -4427 2067
rect -4461 1965 -4427 1999
rect -4461 1897 -4427 1931
rect -4461 1829 -4427 1863
rect -4461 1761 -4427 1795
rect -4461 1693 -4427 1727
rect -4461 1625 -4427 1659
rect -4461 1557 -4427 1591
rect -4461 1489 -4427 1523
rect -4461 1421 -4427 1455
rect -4461 1353 -4427 1387
rect -4461 1285 -4427 1319
rect -4461 1217 -4427 1251
rect -4461 1149 -4427 1183
rect -4461 1081 -4427 1115
rect -4461 1013 -4427 1047
rect -4461 945 -4427 979
rect -4461 877 -4427 911
rect -4461 809 -4427 843
rect -4461 741 -4427 775
rect -4461 673 -4427 707
rect -4461 605 -4427 639
rect -4461 537 -4427 571
rect -4461 469 -4427 503
rect -4461 401 -4427 435
rect -4461 333 -4427 367
rect -4461 265 -4427 299
rect -4461 197 -4427 231
rect -4461 129 -4427 163
rect -4461 61 -4427 95
rect -4461 -7 -4427 27
rect -4461 -75 -4427 -41
rect -4461 -143 -4427 -109
rect -4461 -211 -4427 -177
rect -4461 -279 -4427 -245
rect -4461 -347 -4427 -313
rect -4461 -415 -4427 -381
rect -4461 -483 -4427 -449
rect -4461 -551 -4427 -517
rect -4461 -619 -4427 -585
rect -4461 -687 -4427 -653
rect -4461 -755 -4427 -721
rect -4461 -823 -4427 -789
rect -4461 -891 -4427 -857
rect -4461 -959 -4427 -925
rect -4461 -1027 -4427 -993
rect -4461 -1095 -4427 -1061
rect -4461 -1163 -4427 -1129
rect -4461 -1231 -4427 -1197
rect -4461 -1299 -4427 -1265
rect -4461 -1367 -4427 -1333
rect -4461 -1435 -4427 -1401
rect -4461 -1503 -4427 -1469
rect -4461 -1571 -4427 -1537
rect -4461 -1639 -4427 -1605
rect -4461 -1707 -4427 -1673
rect -4461 -1775 -4427 -1741
rect -4461 -1843 -4427 -1809
rect -4461 -1911 -4427 -1877
rect -4461 -1979 -4427 -1945
rect -4461 -2047 -4427 -2013
rect -4461 -2115 -4427 -2081
rect -4461 -2183 -4427 -2149
rect -4461 -2251 -4427 -2217
rect -4461 -2319 -4427 -2285
rect -4461 -2387 -4427 -2353
rect -4461 -2455 -4427 -2421
rect -4461 -2523 -4427 -2489
rect -4461 -2591 -4427 -2557
rect -4461 -2659 -4427 -2625
rect -4461 -2727 -4427 -2693
rect -4461 -2795 -4427 -2761
rect -4461 -2863 -4427 -2829
rect -4461 -2931 -4427 -2897
rect -4461 -2999 -4427 -2965
rect -4461 -3067 -4427 -3033
rect -4461 -3135 -4427 -3101
rect -4461 -3203 -4427 -3169
rect -4461 -3271 -4427 -3237
rect -4461 -3339 -4427 -3305
rect -4461 -3407 -4427 -3373
rect -4461 -3475 -4427 -3441
rect -4461 -3543 -4427 -3509
rect -4461 -3611 -4427 -3577
rect -4461 -3679 -4427 -3645
rect -4461 -3747 -4427 -3713
rect 2697 6453 2731 6487
rect 2697 6385 2731 6419
rect 2697 6317 2731 6351
rect 2697 6249 2731 6283
rect 2697 6181 2731 6215
rect 2697 6113 2731 6147
rect 2697 6045 2731 6079
rect 2697 5977 2731 6011
rect 2697 5909 2731 5943
rect 2697 5841 2731 5875
rect 2697 5773 2731 5807
rect 2697 5705 2731 5739
rect 2697 5637 2731 5671
rect 2697 5569 2731 5603
rect 2697 5501 2731 5535
rect 2697 5433 2731 5467
rect 2697 5365 2731 5399
rect 2697 5297 2731 5331
rect 2697 5229 2731 5263
rect 2697 5161 2731 5195
rect 2697 5093 2731 5127
rect 2697 5025 2731 5059
rect 2697 4957 2731 4991
rect 2697 4889 2731 4923
rect 2697 4821 2731 4855
rect 2697 4753 2731 4787
rect 2697 4685 2731 4719
rect 2697 4617 2731 4651
rect 2697 4549 2731 4583
rect 2697 4481 2731 4515
rect 2697 4413 2731 4447
rect 2697 4345 2731 4379
rect 2697 4277 2731 4311
rect 2697 4209 2731 4243
rect 2697 4141 2731 4175
rect 2697 4073 2731 4107
rect 2697 4005 2731 4039
rect 2697 3937 2731 3971
rect 2697 3869 2731 3903
rect 2697 3801 2731 3835
rect 2697 3733 2731 3767
rect 2697 3665 2731 3699
rect 2697 3597 2731 3631
rect 2697 3529 2731 3563
rect 2697 3461 2731 3495
rect 2697 3393 2731 3427
rect 2697 3325 2731 3359
rect 2697 3257 2731 3291
rect 2697 3189 2731 3223
rect 2697 3121 2731 3155
rect 2697 3053 2731 3087
rect 2697 2985 2731 3019
rect 2697 2917 2731 2951
rect 2697 2849 2731 2883
rect 2697 2781 2731 2815
rect 2697 2713 2731 2747
rect 2697 2645 2731 2679
rect 2697 2577 2731 2611
rect 2697 2509 2731 2543
rect 2697 2441 2731 2475
rect 2697 2373 2731 2407
rect 2697 2305 2731 2339
rect 2697 2237 2731 2271
rect 2697 2169 2731 2203
rect 2697 2101 2731 2135
rect 2697 2033 2731 2067
rect 2697 1965 2731 1999
rect 2697 1897 2731 1931
rect 2697 1829 2731 1863
rect 2697 1761 2731 1795
rect 2697 1693 2731 1727
rect 2697 1625 2731 1659
rect 2697 1557 2731 1591
rect 2697 1489 2731 1523
rect 2697 1421 2731 1455
rect 2697 1353 2731 1387
rect 2697 1285 2731 1319
rect 2697 1217 2731 1251
rect 2697 1149 2731 1183
rect 2697 1081 2731 1115
rect 2697 1013 2731 1047
rect 2697 945 2731 979
rect 2697 877 2731 911
rect 2697 809 2731 843
rect 2697 741 2731 775
rect 2697 673 2731 707
rect 2697 605 2731 639
rect 2697 537 2731 571
rect 2697 469 2731 503
rect 2697 401 2731 435
rect 2697 333 2731 367
rect 2697 265 2731 299
rect 2697 197 2731 231
rect 2697 129 2731 163
rect 2697 61 2731 95
rect 2697 -7 2731 27
rect 2697 -75 2731 -41
rect 2697 -143 2731 -109
rect 2697 -211 2731 -177
rect 2697 -279 2731 -245
rect 2697 -347 2731 -313
rect 2697 -415 2731 -381
rect 2697 -483 2731 -449
rect 2697 -551 2731 -517
rect 2697 -619 2731 -585
rect 2697 -687 2731 -653
rect 2697 -755 2731 -721
rect 2697 -823 2731 -789
rect 2697 -891 2731 -857
rect 2697 -959 2731 -925
rect 2697 -1027 2731 -993
rect 2697 -1095 2731 -1061
rect 2697 -1163 2731 -1129
rect 2697 -1231 2731 -1197
rect 2697 -1299 2731 -1265
rect 2697 -1367 2731 -1333
rect 2697 -1435 2731 -1401
rect 2697 -1503 2731 -1469
rect 2697 -1571 2731 -1537
rect 2697 -1639 2731 -1605
rect 2697 -1707 2731 -1673
rect 2697 -1775 2731 -1741
rect 2697 -1843 2731 -1809
rect 2697 -1911 2731 -1877
rect 2697 -1979 2731 -1945
rect 2697 -2047 2731 -2013
rect 2697 -2115 2731 -2081
rect 2697 -2183 2731 -2149
rect 2697 -2251 2731 -2217
rect 2697 -2319 2731 -2285
rect 2697 -2387 2731 -2353
rect 2697 -2455 2731 -2421
rect 2697 -2523 2731 -2489
rect 2697 -2591 2731 -2557
rect 2697 -2659 2731 -2625
rect 2697 -2727 2731 -2693
rect 2697 -2795 2731 -2761
rect 2697 -2863 2731 -2829
rect 2697 -2931 2731 -2897
rect 2697 -2999 2731 -2965
rect 2697 -3067 2731 -3033
rect 2697 -3135 2731 -3101
rect 2697 -3203 2731 -3169
rect 2697 -3271 2731 -3237
rect 2697 -3339 2731 -3305
rect 2697 -3407 2731 -3373
rect 2697 -3475 2731 -3441
rect 2697 -3543 2731 -3509
rect 2697 -3611 2731 -3577
rect 2697 -3679 2731 -3645
rect 2697 -3747 2731 -3713
rect -4384 -3815 -4350 -3781
rect -4316 -3815 -4282 -3781
rect -4248 -3815 -4214 -3781
rect -4180 -3815 -4146 -3781
rect -4112 -3815 -4078 -3781
rect -4044 -3815 -4010 -3781
rect -3976 -3815 -3942 -3781
rect -3908 -3815 -3874 -3781
rect -3840 -3815 -3806 -3781
rect -3772 -3815 -3738 -3781
rect -3704 -3815 -3670 -3781
rect -3636 -3815 -3602 -3781
rect -3568 -3815 -3534 -3781
rect -3500 -3815 -3466 -3781
rect -3432 -3815 -3398 -3781
rect -3364 -3815 -3330 -3781
rect -3296 -3815 -3262 -3781
rect -3228 -3815 -3194 -3781
rect -3160 -3815 -3126 -3781
rect -3092 -3815 -3058 -3781
rect -3024 -3815 -2990 -3781
rect -2956 -3815 -2922 -3781
rect -2888 -3815 -2854 -3781
rect -2820 -3815 -2786 -3781
rect -2752 -3815 -2718 -3781
rect -2684 -3815 -2650 -3781
rect -2616 -3815 -2582 -3781
rect -2548 -3815 -2514 -3781
rect -2480 -3815 -2446 -3781
rect -2412 -3815 -2378 -3781
rect -2344 -3815 -2310 -3781
rect -2276 -3815 -2242 -3781
rect -2208 -3815 -2174 -3781
rect -2140 -3815 -2106 -3781
rect -2072 -3815 -2038 -3781
rect -2004 -3815 -1970 -3781
rect -1936 -3815 -1902 -3781
rect -1868 -3815 -1834 -3781
rect -1800 -3815 -1766 -3781
rect -1732 -3815 -1698 -3781
rect -1664 -3815 -1630 -3781
rect -1596 -3815 -1562 -3781
rect -1528 -3815 -1494 -3781
rect -1460 -3815 -1426 -3781
rect -1392 -3815 -1358 -3781
rect -1324 -3815 -1290 -3781
rect -1256 -3815 -1222 -3781
rect -1188 -3815 -1154 -3781
rect -1120 -3815 -1086 -3781
rect -1052 -3815 -1018 -3781
rect -984 -3815 -950 -3781
rect -916 -3815 -882 -3781
rect -848 -3815 -814 -3781
rect -780 -3815 -746 -3781
rect -712 -3815 -678 -3781
rect -644 -3815 -610 -3781
rect -576 -3815 -542 -3781
rect -508 -3815 -474 -3781
rect -440 -3815 -406 -3781
rect -372 -3815 -338 -3781
rect -304 -3815 -270 -3781
rect -236 -3815 -202 -3781
rect -168 -3815 -134 -3781
rect -100 -3815 -66 -3781
rect -32 -3815 2 -3781
rect 36 -3815 70 -3781
rect 104 -3815 138 -3781
rect 172 -3815 206 -3781
rect 240 -3815 274 -3781
rect 308 -3815 342 -3781
rect 376 -3815 410 -3781
rect 444 -3815 478 -3781
rect 512 -3815 546 -3781
rect 580 -3815 614 -3781
rect 648 -3815 682 -3781
rect 716 -3815 750 -3781
rect 784 -3815 818 -3781
rect 852 -3815 886 -3781
rect 920 -3815 954 -3781
rect 988 -3815 1022 -3781
rect 1056 -3815 1090 -3781
rect 1124 -3815 1158 -3781
rect 1192 -3815 1226 -3781
rect 1260 -3815 1294 -3781
rect 1328 -3815 1362 -3781
rect 1396 -3815 1430 -3781
rect 1464 -3815 1498 -3781
rect 1532 -3815 1566 -3781
rect 1600 -3815 1634 -3781
rect 1668 -3815 1702 -3781
rect 1736 -3815 1770 -3781
rect 1804 -3815 1838 -3781
rect 1872 -3815 1906 -3781
rect 1940 -3815 1974 -3781
rect 2008 -3815 2042 -3781
rect 2076 -3815 2110 -3781
rect 2144 -3815 2178 -3781
rect 2212 -3815 2246 -3781
rect 2280 -3815 2314 -3781
rect 2348 -3815 2382 -3781
rect 2416 -3815 2450 -3781
rect 2484 -3815 2518 -3781
rect 2552 -3815 2586 -3781
rect 2620 -3815 2654 -3781
<< locali >>
rect -4461 6521 -4384 6555
rect -4350 6521 -4316 6555
rect -4282 6521 -4248 6555
rect -4214 6521 -4180 6555
rect -4146 6521 -4112 6555
rect -4078 6521 -4044 6555
rect -4010 6521 -3976 6555
rect -3942 6521 -3908 6555
rect -3874 6521 -3840 6555
rect -3806 6521 -3772 6555
rect -3738 6521 -3704 6555
rect -3670 6521 -3636 6555
rect -3602 6521 -3568 6555
rect -3534 6521 -3500 6555
rect -3466 6521 -3432 6555
rect -3398 6521 -3364 6555
rect -3330 6521 -3296 6555
rect -3262 6521 -3228 6555
rect -3194 6521 -3160 6555
rect -3126 6521 -3092 6555
rect -3058 6521 -3024 6555
rect -2990 6521 -2956 6555
rect -2922 6521 -2888 6555
rect -2854 6521 -2820 6555
rect -2786 6521 -2752 6555
rect -2718 6521 -2684 6555
rect -2650 6521 -2616 6555
rect -2582 6521 -2548 6555
rect -2514 6521 -2480 6555
rect -2446 6521 -2412 6555
rect -2378 6521 -2344 6555
rect -2310 6521 -2276 6555
rect -2242 6521 -2208 6555
rect -2174 6521 -2140 6555
rect -2106 6521 -2072 6555
rect -2038 6521 -2004 6555
rect -1970 6521 -1936 6555
rect -1902 6521 -1868 6555
rect -1834 6521 -1800 6555
rect -1766 6521 -1732 6555
rect -1698 6521 -1664 6555
rect -1630 6521 -1596 6555
rect -1562 6521 -1528 6555
rect -1494 6521 -1460 6555
rect -1426 6521 -1392 6555
rect -1358 6521 -1324 6555
rect -1290 6521 -1256 6555
rect -1222 6521 -1188 6555
rect -1154 6521 -1120 6555
rect -1086 6521 -1052 6555
rect -1018 6521 -984 6555
rect -950 6521 -916 6555
rect -882 6521 -848 6555
rect -814 6521 -780 6555
rect -746 6521 -712 6555
rect -678 6521 -644 6555
rect -610 6521 -576 6555
rect -542 6521 -508 6555
rect -474 6521 -440 6555
rect -406 6521 -372 6555
rect -338 6521 -304 6555
rect -270 6521 -236 6555
rect -202 6521 -168 6555
rect -134 6521 -100 6555
rect -66 6521 -32 6555
rect 2 6521 36 6555
rect 70 6521 104 6555
rect 138 6521 172 6555
rect 206 6521 240 6555
rect 274 6521 308 6555
rect 342 6521 376 6555
rect 410 6521 444 6555
rect 478 6521 512 6555
rect 546 6521 580 6555
rect 614 6521 648 6555
rect 682 6521 716 6555
rect 750 6521 784 6555
rect 818 6521 852 6555
rect 886 6521 920 6555
rect 954 6521 988 6555
rect 1022 6521 1056 6555
rect 1090 6521 1124 6555
rect 1158 6521 1192 6555
rect 1226 6521 1260 6555
rect 1294 6521 1328 6555
rect 1362 6521 1396 6555
rect 1430 6521 1464 6555
rect 1498 6521 1532 6555
rect 1566 6521 1600 6555
rect 1634 6521 1668 6555
rect 1702 6521 1736 6555
rect 1770 6521 1804 6555
rect 1838 6521 1872 6555
rect 1906 6521 1940 6555
rect 1974 6521 2008 6555
rect 2042 6521 2076 6555
rect 2110 6521 2144 6555
rect 2178 6521 2212 6555
rect 2246 6521 2280 6555
rect 2314 6521 2348 6555
rect 2382 6521 2416 6555
rect 2450 6521 2484 6555
rect 2518 6521 2552 6555
rect 2586 6521 2620 6555
rect 2654 6521 2731 6555
rect -4461 6487 2731 6521
rect -4427 6470 2697 6487
rect -4427 6453 -4317 6470
rect -4461 6419 -4317 6453
rect -4427 6385 -4317 6419
rect -4461 6364 -4317 6385
rect 2629 6453 2697 6470
rect 2629 6419 2731 6453
rect 2629 6385 2697 6419
rect 2629 6364 2731 6385
rect -4461 6351 2731 6364
rect -4427 6317 2697 6351
rect -4461 6296 2731 6317
rect -4461 6283 -4318 6296
rect -4427 6262 -4318 6283
rect -4284 6283 2731 6296
rect -4284 6262 2697 6283
rect -4427 6252 2697 6262
rect -4427 6249 -4147 6252
rect -4461 6224 -4147 6249
rect -4461 6215 -4318 6224
rect -4427 6190 -4318 6215
rect -4284 6190 -4147 6224
rect -4427 6181 -4147 6190
rect -4461 6152 -4147 6181
rect -4461 6147 -4318 6152
rect -4427 6118 -4318 6147
rect -4284 6118 -4147 6152
rect -4427 6113 -4147 6118
rect -4461 6080 -4147 6113
rect -4461 6079 -4318 6080
rect -4427 6046 -4318 6079
rect -4284 6046 -4147 6080
rect -4427 6045 -4147 6046
rect -4461 6011 -4147 6045
rect -4427 6008 -4147 6011
rect -4427 5977 -4318 6008
rect -4461 5974 -4318 5977
rect -4284 5974 -4147 6008
rect -4461 5943 -4147 5974
rect -4427 5936 -4147 5943
rect -4427 5909 -4318 5936
rect -4461 5902 -4318 5909
rect -4284 5902 -4147 5936
rect -4461 5875 -4147 5902
rect -4427 5864 -4147 5875
rect -4427 5841 -4318 5864
rect -4461 5830 -4318 5841
rect -4284 5830 -4147 5864
rect -4461 5807 -4147 5830
rect -4427 5792 -4147 5807
rect -4427 5773 -4318 5792
rect -4461 5758 -4318 5773
rect -4284 5758 -4147 5792
rect -4461 5739 -4147 5758
rect -4427 5720 -4147 5739
rect -4427 5705 -4318 5720
rect -4461 5686 -4318 5705
rect -4284 5686 -4147 5720
rect -4461 5671 -4147 5686
rect -4427 5648 -4147 5671
rect -4427 5637 -4318 5648
rect -4461 5614 -4318 5637
rect -4284 5614 -4147 5648
rect -4461 5603 -4147 5614
rect -4427 5576 -4147 5603
rect -4427 5569 -4318 5576
rect -4461 5542 -4318 5569
rect -4284 5542 -4147 5576
rect -4461 5535 -4147 5542
rect -4427 5504 -4147 5535
rect -4427 5501 -4318 5504
rect -4461 5470 -4318 5501
rect -4284 5470 -4147 5504
rect -4461 5467 -4147 5470
rect -4427 5433 -4147 5467
rect -4461 5432 -4147 5433
rect -4461 5399 -4318 5432
rect -4427 5398 -4318 5399
rect -4284 5398 -4147 5432
rect -4427 5365 -4147 5398
rect -4461 5360 -4147 5365
rect -4461 5331 -4318 5360
rect -4427 5326 -4318 5331
rect -4284 5326 -4147 5360
rect -4427 5297 -4147 5326
rect -4461 5288 -4147 5297
rect -4461 5263 -4318 5288
rect -4427 5254 -4318 5263
rect -4284 5254 -4147 5288
rect -4427 5229 -4147 5254
rect -4461 5216 -4147 5229
rect -4461 5195 -4318 5216
rect -4427 5182 -4318 5195
rect -4284 5182 -4147 5216
rect -4427 5161 -4147 5182
rect -4461 5144 -4147 5161
rect -4461 5127 -4318 5144
rect -4427 5110 -4318 5127
rect -4284 5110 -4147 5144
rect -4427 5093 -4147 5110
rect -4461 5072 -4147 5093
rect -4461 5059 -4318 5072
rect -4427 5038 -4318 5059
rect -4284 5038 -4147 5072
rect -4427 5025 -4147 5038
rect -4461 5000 -4147 5025
rect -4461 4991 -4318 5000
rect -4427 4966 -4318 4991
rect -4284 4966 -4147 5000
rect -4427 4957 -4147 4966
rect -4461 4928 -4147 4957
rect -4461 4923 -4318 4928
rect -4427 4894 -4318 4923
rect -4284 4894 -4147 4928
rect -4427 4889 -4147 4894
rect -4461 4856 -4147 4889
rect -4461 4855 -4318 4856
rect -4427 4822 -4318 4855
rect -4284 4822 -4147 4856
rect -4427 4821 -4147 4822
rect -4461 4787 -4147 4821
rect -4427 4784 -4147 4787
rect -4427 4753 -4318 4784
rect -4461 4750 -4318 4753
rect -4284 4750 -4147 4784
rect -4461 4719 -4147 4750
rect -4427 4712 -4147 4719
rect -4427 4685 -4318 4712
rect -4461 4678 -4318 4685
rect -4284 4678 -4147 4712
rect -4461 4651 -4147 4678
rect -4427 4640 -4147 4651
rect -4427 4617 -4318 4640
rect -4461 4606 -4318 4617
rect -4284 4606 -4147 4640
rect -4461 4583 -4147 4606
rect -4427 4568 -4147 4583
rect -4427 4549 -4318 4568
rect -4461 4534 -4318 4549
rect -4284 4534 -4147 4568
rect -4461 4515 -4147 4534
rect -4427 4496 -4147 4515
rect -4427 4481 -4318 4496
rect -4461 4462 -4318 4481
rect -4284 4462 -4147 4496
rect -4461 4447 -4147 4462
rect -4427 4424 -4147 4447
rect -4427 4413 -4318 4424
rect -4461 4390 -4318 4413
rect -4284 4390 -4147 4424
rect -4461 4379 -4147 4390
rect -4427 4352 -4147 4379
rect -4427 4345 -4318 4352
rect -4461 4318 -4318 4345
rect -4284 4318 -4147 4352
rect -4461 4311 -4147 4318
rect -4427 4280 -4147 4311
rect -4427 4277 -4318 4280
rect -4461 4246 -4318 4277
rect -4284 4246 -4147 4280
rect -4461 4243 -4147 4246
rect -4427 4209 -4147 4243
rect -4461 4208 -4147 4209
rect -4461 4175 -4318 4208
rect -4427 4174 -4318 4175
rect -4284 4174 -4147 4208
rect -4427 4141 -4147 4174
rect -4461 4107 -4147 4141
rect -4427 4073 -4147 4107
rect -4461 4039 -4147 4073
rect -4427 4005 -4147 4039
rect -4461 3971 -4147 4005
rect -4427 3937 -4147 3971
rect -4461 3929 -4147 3937
rect 2432 6249 2697 6252
rect 2432 6215 2731 6249
rect 2432 6181 2697 6215
rect 2432 6147 2731 6181
rect 2432 6113 2697 6147
rect 2432 6079 2731 6113
rect 2432 6045 2697 6079
rect 2432 6011 2731 6045
rect 2432 5977 2697 6011
rect 2432 5943 2731 5977
rect 2432 5909 2697 5943
rect 2432 5875 2731 5909
rect 2432 5841 2697 5875
rect 2432 5807 2731 5841
rect 2432 5773 2697 5807
rect 2432 5739 2731 5773
rect 2432 5705 2697 5739
rect 2432 5671 2731 5705
rect 2432 5637 2697 5671
rect 2432 5603 2731 5637
rect 2432 5569 2697 5603
rect 2432 5535 2731 5569
rect 2432 5501 2697 5535
rect 2432 5467 2731 5501
rect 2432 5433 2697 5467
rect 2432 5399 2731 5433
rect 2432 5365 2697 5399
rect 2432 5331 2731 5365
rect 2432 5297 2697 5331
rect 2432 5263 2731 5297
rect 2432 5229 2697 5263
rect 2432 5195 2731 5229
rect 2432 5161 2697 5195
rect 2432 5127 2731 5161
rect 2432 5093 2697 5127
rect 2432 5059 2731 5093
rect 2432 5025 2697 5059
rect 2432 4991 2731 5025
rect 2432 4957 2697 4991
rect 2432 4923 2731 4957
rect 2432 4889 2697 4923
rect 2432 4855 2731 4889
rect 2432 4821 2697 4855
rect 2432 4787 2731 4821
rect 2432 4753 2697 4787
rect 2432 4719 2731 4753
rect 2432 4685 2697 4719
rect 2432 4651 2731 4685
rect 2432 4617 2697 4651
rect 2432 4583 2731 4617
rect 2432 4549 2697 4583
rect 2432 4515 2731 4549
rect 2432 4481 2697 4515
rect 2432 4447 2731 4481
rect 2432 4413 2697 4447
rect 2432 4379 2731 4413
rect 2432 4345 2697 4379
rect 2432 4311 2731 4345
rect 2432 4277 2697 4311
rect 2432 4243 2731 4277
rect 2432 4209 2697 4243
rect 2432 4175 2731 4209
rect 2432 4141 2697 4175
rect 2432 4107 2731 4141
rect 2432 4073 2697 4107
rect 2432 4039 2731 4073
rect 2432 4005 2697 4039
rect 2432 3971 2731 4005
rect 2432 3937 2697 3971
rect 2432 3929 2731 3937
rect -4461 3926 2731 3929
rect -4461 3903 -4148 3926
rect -4427 3892 -4148 3903
rect -4114 3892 -4076 3926
rect -4042 3892 -4004 3926
rect -3970 3892 -3932 3926
rect -3898 3892 -3860 3926
rect -3826 3892 -3788 3926
rect -3754 3892 -3716 3926
rect -3682 3892 -3644 3926
rect -3610 3892 -3572 3926
rect -3538 3892 -3500 3926
rect -3466 3892 -3428 3926
rect -3394 3892 -3356 3926
rect -3322 3892 -3284 3926
rect -3250 3892 -3212 3926
rect -3178 3892 -3140 3926
rect -3106 3892 -3068 3926
rect -3034 3892 -2996 3926
rect -2962 3892 -2924 3926
rect -2890 3892 -2852 3926
rect -2818 3892 -2780 3926
rect -2746 3892 -2708 3926
rect -2674 3892 -2636 3926
rect -2602 3892 -2564 3926
rect -2530 3892 -2492 3926
rect -2458 3892 -2420 3926
rect -2386 3892 -2348 3926
rect -2314 3892 -2276 3926
rect -2242 3892 -2204 3926
rect -2170 3892 -2132 3926
rect -2098 3892 -2060 3926
rect -2026 3892 -1988 3926
rect -1954 3892 -1916 3926
rect -1882 3892 -1844 3926
rect -1810 3892 -1772 3926
rect -1738 3892 -1700 3926
rect -1666 3892 -1628 3926
rect -1594 3892 -1556 3926
rect -1522 3892 -1484 3926
rect -1450 3892 -1412 3926
rect -1378 3892 -1340 3926
rect -1306 3892 -1268 3926
rect -1234 3892 -1196 3926
rect -1162 3892 -1124 3926
rect -1090 3892 -1052 3926
rect -1018 3892 -980 3926
rect -946 3892 -908 3926
rect -874 3892 -836 3926
rect -802 3892 -764 3926
rect -730 3892 -692 3926
rect -658 3892 -620 3926
rect -586 3892 -548 3926
rect -514 3892 -476 3926
rect -442 3892 -404 3926
rect -370 3892 -332 3926
rect -298 3892 -260 3926
rect -226 3892 -188 3926
rect -154 3892 -116 3926
rect -82 3892 -44 3926
rect -10 3892 28 3926
rect 62 3892 100 3926
rect 134 3892 172 3926
rect 206 3892 244 3926
rect 278 3892 316 3926
rect 350 3892 388 3926
rect 422 3892 460 3926
rect 494 3892 532 3926
rect 566 3892 604 3926
rect 638 3892 676 3926
rect 710 3892 748 3926
rect 782 3892 820 3926
rect 854 3892 892 3926
rect 926 3892 964 3926
rect 998 3892 1036 3926
rect 1070 3892 1108 3926
rect 1142 3892 1180 3926
rect 1214 3892 1252 3926
rect 1286 3892 1324 3926
rect 1358 3892 1396 3926
rect 1430 3892 1468 3926
rect 1502 3892 1540 3926
rect 1574 3892 1612 3926
rect 1646 3892 1684 3926
rect 1718 3892 1756 3926
rect 1790 3892 1828 3926
rect 1862 3892 1900 3926
rect 1934 3892 1972 3926
rect 2006 3892 2044 3926
rect 2078 3892 2116 3926
rect 2150 3892 2188 3926
rect 2222 3892 2260 3926
rect 2294 3892 2332 3926
rect 2366 3892 2404 3926
rect 2438 3903 2731 3926
rect 2438 3892 2697 3903
rect -4427 3889 2697 3892
rect -4427 3869 -4147 3889
rect -4461 3835 -4147 3869
rect -4427 3801 -4147 3835
rect -4461 3767 -4147 3801
rect -4427 3733 -4147 3767
rect -4461 3699 -4147 3733
rect -4427 3665 -4147 3699
rect -4461 3631 -4147 3665
rect -4427 3597 -4147 3631
rect -4461 3563 -4147 3597
rect -4427 3529 -4147 3563
rect -4461 3495 -4147 3529
rect -4427 3461 -4147 3495
rect -4461 3427 -4147 3461
rect -4427 3393 -4147 3427
rect -4461 3359 -4147 3393
rect -4427 3325 -4147 3359
rect -4461 3291 -4147 3325
rect -4427 3257 -4147 3291
rect -4461 3223 -4147 3257
rect -4427 3189 -4147 3223
rect -4461 3155 -4147 3189
rect -4427 3121 -4147 3155
rect -4461 3087 -4147 3121
rect -4427 3053 -4147 3087
rect -4461 3019 -4147 3053
rect -4427 2985 -4147 3019
rect -4461 2951 -4147 2985
rect -4427 2917 -4147 2951
rect -4461 2883 -4147 2917
rect -4427 2849 -4147 2883
rect -4461 2815 -4147 2849
rect -4427 2781 -4147 2815
rect -4461 2747 -4147 2781
rect -4427 2713 -4147 2747
rect -4461 2679 -4147 2713
rect -4427 2645 -4147 2679
rect -4461 2611 -4147 2645
rect -4427 2577 -4147 2611
rect -4461 2543 -4147 2577
rect -4427 2509 -4147 2543
rect -4461 2475 -4147 2509
rect -4427 2441 -4147 2475
rect -4461 2407 -4147 2441
rect -4427 2373 -4147 2407
rect -4461 2339 -4147 2373
rect -4427 2305 -4147 2339
rect -4461 2271 -4147 2305
rect -4427 2237 -4147 2271
rect -4461 2203 -4147 2237
rect -4427 2169 -4147 2203
rect -4461 2135 -4147 2169
rect -4427 2101 -4147 2135
rect -4461 2067 -4147 2101
rect -4427 2033 -4147 2067
rect -4461 1999 -4147 2033
rect -4427 1965 -4147 1999
rect -4461 1931 -4147 1965
rect -4427 1897 -4147 1931
rect -4461 1863 -4147 1897
rect -4427 1829 -4147 1863
rect -4461 1795 -4147 1829
rect -4427 1761 -4147 1795
rect -4461 1727 -4147 1761
rect -4427 1693 -4147 1727
rect -4461 1659 -4147 1693
rect -4427 1625 -4147 1659
rect -4461 1591 -4147 1625
rect -4427 1567 -4147 1591
rect 2432 3869 2697 3889
rect 2432 3835 2731 3869
rect 2432 3801 2697 3835
rect 2432 3767 2731 3801
rect 2432 3733 2697 3767
rect 2432 3699 2731 3733
rect 2432 3665 2697 3699
rect 2432 3631 2731 3665
rect 2432 3597 2697 3631
rect 2432 3563 2731 3597
rect 2432 3529 2697 3563
rect 2432 3495 2731 3529
rect 2432 3461 2697 3495
rect 2432 3427 2731 3461
rect 2432 3393 2697 3427
rect 2432 3359 2731 3393
rect 2432 3325 2697 3359
rect 2432 3291 2731 3325
rect 2432 3257 2697 3291
rect 2432 3223 2731 3257
rect 2432 3189 2697 3223
rect 2432 3155 2731 3189
rect 2432 3121 2697 3155
rect 2432 3087 2731 3121
rect 2432 3053 2697 3087
rect 2432 3019 2731 3053
rect 2432 2985 2697 3019
rect 2432 2951 2731 2985
rect 2432 2917 2697 2951
rect 2432 2883 2731 2917
rect 2432 2849 2697 2883
rect 2432 2815 2731 2849
rect 2432 2781 2697 2815
rect 2432 2747 2731 2781
rect 2432 2713 2697 2747
rect 2432 2679 2731 2713
rect 2432 2645 2697 2679
rect 2432 2611 2731 2645
rect 2432 2577 2697 2611
rect 2432 2543 2731 2577
rect 2432 2509 2697 2543
rect 2432 2475 2731 2509
rect 2432 2441 2697 2475
rect 2432 2407 2731 2441
rect 2432 2373 2697 2407
rect 2432 2339 2731 2373
rect 2432 2305 2697 2339
rect 2432 2271 2731 2305
rect 2432 2237 2697 2271
rect 2432 2203 2731 2237
rect 2432 2169 2697 2203
rect 2432 2135 2731 2169
rect 2432 2101 2697 2135
rect 2432 2067 2731 2101
rect 2432 2033 2697 2067
rect 2432 1999 2731 2033
rect 2432 1965 2697 1999
rect 2432 1931 2731 1965
rect 2432 1897 2697 1931
rect 2432 1863 2731 1897
rect 2432 1829 2697 1863
rect 2432 1795 2731 1829
rect 2432 1761 2697 1795
rect 2432 1727 2731 1761
rect 2432 1693 2697 1727
rect 2432 1659 2731 1693
rect 2432 1625 2697 1659
rect 2432 1591 2731 1625
rect 2432 1567 2697 1591
rect -4427 1557 2697 1567
rect -4461 1523 2731 1557
rect -4427 1489 2697 1523
rect -4461 1455 2731 1489
rect -4427 1421 2697 1455
rect -4461 1401 2731 1421
rect -4461 1400 2148 1401
rect -4461 1399 1404 1400
rect -4461 1387 -4035 1399
rect -4427 1353 -4035 1387
rect -4461 1319 -4035 1353
rect -4427 1285 -4035 1319
rect -4461 1251 -4035 1285
rect -4427 1221 -4035 1251
rect -3857 1381 1404 1399
rect -3857 1221 -3397 1381
rect -4427 1217 -3397 1221
rect -4461 1183 -3397 1217
rect -4427 1179 -3397 1183
rect -4427 1149 -4342 1179
rect -4461 1115 -4342 1149
rect -4427 1081 -4342 1115
rect -4461 1047 -4342 1081
rect -4427 1013 -4342 1047
rect -4461 979 -4342 1013
rect -4427 945 -4342 979
rect -4461 929 -4342 945
rect -4164 965 -3397 1179
rect -4164 929 -4140 965
rect -4461 911 -4140 929
rect -4427 877 -4140 911
rect -4461 843 -4140 877
rect -4427 809 -4140 843
rect -4461 775 -4140 809
rect -4427 741 -4140 775
rect -4461 707 -4140 741
rect -4427 673 -4140 707
rect -4461 639 -4140 673
rect -4427 605 -4140 639
rect -4461 571 -4140 605
rect -4427 537 -4140 571
rect -4461 503 -4140 537
rect -4427 469 -4140 503
rect -4461 435 -4140 469
rect -4427 401 -4140 435
rect -4461 367 -4140 401
rect -4427 333 -4140 367
rect -4461 299 -4140 333
rect -4427 265 -4140 299
rect -4461 231 -4140 265
rect -4427 197 -4140 231
rect -4461 164 -4140 197
rect -4060 649 -3579 889
rect -4060 354 -3950 649
rect -3660 354 -3579 649
rect -3495 555 -3397 965
rect -3291 1366 1404 1381
rect -3291 1260 -3193 1366
rect 1305 1260 1404 1366
rect -3291 959 1404 1260
rect -3291 555 -3196 959
rect -3495 420 -3196 555
rect 1313 502 1404 959
rect 1510 1223 2148 1400
rect 2326 1387 2731 1401
rect 2326 1353 2697 1387
rect 2326 1319 2731 1353
rect 2326 1285 2697 1319
rect 2326 1251 2731 1285
rect 2326 1223 2697 1251
rect 1510 1217 2697 1223
rect 1510 1183 2731 1217
rect 1510 1149 2697 1183
rect 1510 1115 2731 1149
rect 1510 1081 2697 1115
rect 1510 1047 2731 1081
rect 1510 1013 2697 1047
rect 1510 979 2731 1013
rect 1510 954 2697 979
rect 1510 502 1610 954
rect 1313 420 1610 502
rect -3495 363 1610 420
rect 2374 945 2697 954
rect 2374 911 2731 945
rect 2374 877 2697 911
rect 2374 843 2731 877
rect 2374 809 2697 843
rect 2374 775 2731 809
rect 2374 741 2697 775
rect 2374 707 2731 741
rect 2374 673 2697 707
rect 2374 639 2731 673
rect 2374 605 2697 639
rect 2374 571 2731 605
rect 2374 537 2697 571
rect 2374 503 2731 537
rect 2374 469 2697 503
rect 2374 435 2731 469
rect 2374 401 2697 435
rect 2374 367 2731 401
rect -4060 197 -3579 354
rect 2374 333 2697 367
rect 2374 299 2731 333
rect 2374 265 2697 299
rect 2374 231 2731 265
rect 2374 197 2697 231
rect -4461 163 -4296 164
rect -4427 129 -4296 163
rect -4461 95 -4296 129
rect -4427 61 -4296 95
rect -4060 152 2291 197
rect 2374 188 2731 197
rect -4060 62 -3306 152
rect -4461 27 -4296 61
rect -4427 -7 -4296 27
rect -4461 -41 -4296 -7
rect -4427 -75 -4296 -41
rect -4461 -109 -4296 -75
rect -4427 -143 -4296 -109
rect -4461 -177 -4296 -143
rect -4427 -211 -4296 -177
rect -4461 -245 -4296 -211
rect -4427 -279 -4296 -245
rect -4184 50 -3306 62
rect -4184 15 -3931 50
rect -4184 -246 -4105 15
rect -4461 -313 -4296 -279
rect -4427 -347 -4296 -313
rect -4461 -381 -4296 -347
rect -4427 -415 -4296 -381
rect -4461 -449 -4296 -415
rect -4183 -440 -4105 -246
rect -4427 -483 -4296 -449
rect -4461 -517 -4296 -483
rect -4427 -551 -4296 -517
rect -4461 -585 -4296 -551
rect -4427 -619 -4296 -585
rect -4461 -653 -4296 -619
rect -4427 -667 -4296 -653
rect -4427 -687 -4382 -667
rect -4461 -701 -4382 -687
rect -4348 -701 -4296 -667
rect -4186 -523 -4105 -440
rect -3999 -239 -3931 15
rect -3658 15 -3306 50
rect -3658 -239 -3509 15
rect -3999 -451 -3509 -239
rect -3403 -440 -3306 15
rect 1918 109 2291 152
rect 2561 163 2731 188
rect 2561 129 2697 163
rect 1918 -440 2440 109
rect -3403 -451 2440 -440
rect -3999 -518 2440 -451
rect 2561 95 2731 129
rect 2561 61 2697 95
rect 2561 27 2731 61
rect 2561 -7 2697 27
rect 2561 -41 2731 -7
rect 2561 -75 2697 -41
rect 2561 -109 2731 -75
rect 2561 -143 2697 -109
rect 2561 -177 2731 -143
rect 2561 -211 2697 -177
rect 2561 -245 2731 -211
rect 2561 -279 2697 -245
rect 2561 -313 2731 -279
rect 2561 -347 2697 -313
rect 2561 -381 2731 -347
rect 2561 -415 2697 -381
rect 2561 -449 2731 -415
rect 2561 -483 2697 -449
rect 2561 -517 2731 -483
rect -3999 -523 2439 -518
rect -4186 -583 2439 -523
rect -4186 -617 -3652 -583
rect -3618 -617 -3580 -583
rect -3546 -617 -3508 -583
rect -3474 -617 -3436 -583
rect -3402 -617 -3364 -583
rect -3330 -617 -3292 -583
rect -3258 -617 -3220 -583
rect -3186 -617 -3148 -583
rect -3114 -617 -3076 -583
rect -3042 -617 -3004 -583
rect -2970 -617 -2932 -583
rect -2898 -617 -2860 -583
rect -2826 -617 -2788 -583
rect -2754 -617 -2716 -583
rect -2682 -617 -2644 -583
rect -2610 -617 -2572 -583
rect -2538 -617 -2500 -583
rect -2466 -617 -2428 -583
rect -2394 -617 -2356 -583
rect -2322 -617 -2284 -583
rect -2250 -617 -2212 -583
rect -2178 -617 -2140 -583
rect -2106 -617 -2068 -583
rect -2034 -617 -1996 -583
rect -1962 -617 -1924 -583
rect -1890 -617 -1852 -583
rect -1818 -617 -1780 -583
rect -1746 -617 -1708 -583
rect -1674 -617 -1636 -583
rect -1602 -617 -1564 -583
rect -1530 -617 -1492 -583
rect -1458 -617 -1420 -583
rect -1386 -617 -1348 -583
rect -1314 -617 -1276 -583
rect -1242 -617 -1204 -583
rect -1170 -617 -1132 -583
rect -1098 -617 -1060 -583
rect -1026 -617 -988 -583
rect -954 -617 -916 -583
rect -882 -617 -844 -583
rect -810 -617 -772 -583
rect -738 -617 -700 -583
rect -666 -617 -628 -583
rect -594 -617 -556 -583
rect -522 -617 -484 -583
rect -450 -617 -412 -583
rect -378 -617 -340 -583
rect -306 -617 -268 -583
rect -234 -617 -196 -583
rect -162 -617 -124 -583
rect -90 -617 -52 -583
rect -18 -617 20 -583
rect 54 -617 92 -583
rect 126 -617 164 -583
rect 198 -617 236 -583
rect 270 -617 308 -583
rect 342 -617 380 -583
rect 414 -617 452 -583
rect 486 -617 524 -583
rect 558 -617 596 -583
rect 630 -617 668 -583
rect 702 -617 740 -583
rect 774 -617 812 -583
rect 846 -617 884 -583
rect 918 -617 956 -583
rect 990 -617 1028 -583
rect 1062 -617 1100 -583
rect 1134 -617 1172 -583
rect 1206 -617 1244 -583
rect 1278 -617 1316 -583
rect 1350 -617 1388 -583
rect 1422 -617 1460 -583
rect 1494 -617 1532 -583
rect 1566 -617 1604 -583
rect 1638 -617 1676 -583
rect 1710 -617 1748 -583
rect 1782 -617 1820 -583
rect 1854 -617 1892 -583
rect 1926 -617 1964 -583
rect 1998 -617 2036 -583
rect 2070 -617 2108 -583
rect 2142 -617 2180 -583
rect 2214 -617 2439 -583
rect -4186 -680 2439 -617
rect 2561 -551 2697 -517
rect 2561 -585 2731 -551
rect 2561 -619 2697 -585
rect 2561 -653 2731 -619
rect -4461 -721 -4296 -701
rect -4427 -739 -4296 -721
rect -4427 -755 -4382 -739
rect -4461 -773 -4382 -755
rect -4348 -773 -4296 -739
rect -4461 -789 -4296 -773
rect -4427 -811 -4296 -789
rect -4427 -823 -4382 -811
rect -4461 -845 -4382 -823
rect -4348 -845 -4296 -811
rect -4461 -857 -4296 -845
rect -4427 -883 -4296 -857
rect -4427 -891 -4382 -883
rect -4461 -917 -4382 -891
rect -4348 -917 -4296 -883
rect -4461 -925 -4296 -917
rect -4427 -955 -4296 -925
rect -4427 -959 -4382 -955
rect -4461 -989 -4382 -959
rect -4348 -989 -4296 -955
rect -4461 -993 -4296 -989
rect -4427 -1027 -4296 -993
rect -4461 -1061 -4382 -1027
rect -4348 -1061 -4296 -1027
rect -4427 -1095 -4296 -1061
rect -4461 -1099 -4296 -1095
rect -4461 -1129 -4382 -1099
rect -4427 -1133 -4382 -1129
rect -4348 -1133 -4296 -1099
rect -4427 -1163 -4296 -1133
rect -4461 -1171 -4296 -1163
rect -4461 -1197 -4382 -1171
rect -4427 -1205 -4382 -1197
rect -4348 -1205 -4296 -1171
rect -4427 -1231 -4296 -1205
rect -4461 -1243 -4296 -1231
rect -4461 -1265 -4382 -1243
rect -4427 -1277 -4382 -1265
rect -4348 -1277 -4296 -1243
rect -4427 -1299 -4296 -1277
rect -4461 -1315 -4296 -1299
rect -4461 -1333 -4382 -1315
rect -4427 -1349 -4382 -1333
rect -4348 -1349 -4296 -1315
rect -4427 -1367 -4296 -1349
rect -4461 -1387 -4296 -1367
rect -4461 -1401 -4382 -1387
rect -4427 -1421 -4382 -1401
rect -4348 -1421 -4296 -1387
rect -4427 -1435 -4296 -1421
rect -4461 -1459 -4296 -1435
rect -4461 -1469 -4382 -1459
rect -4427 -1493 -4382 -1469
rect -4348 -1493 -4296 -1459
rect -4427 -1503 -4296 -1493
rect -4461 -1531 -4296 -1503
rect -4461 -1537 -4382 -1531
rect -4427 -1565 -4382 -1537
rect -4348 -1565 -4296 -1531
rect -4427 -1571 -4296 -1565
rect -4461 -1603 -4296 -1571
rect -4461 -1605 -4382 -1603
rect -4427 -1637 -4382 -1605
rect -4348 -1637 -4296 -1603
rect -4427 -1639 -4296 -1637
rect -4461 -1673 -4296 -1639
rect -4427 -1675 -4296 -1673
rect -4427 -1707 -4382 -1675
rect -4461 -1709 -4382 -1707
rect -4348 -1709 -4296 -1675
rect -4461 -1741 -4296 -1709
rect -4427 -1747 -4296 -1741
rect -4427 -1775 -4382 -1747
rect -4461 -1781 -4382 -1775
rect -4348 -1781 -4296 -1747
rect -4461 -1809 -4296 -1781
rect -4427 -1819 -4296 -1809
rect -4427 -1843 -4382 -1819
rect -4461 -1853 -4382 -1843
rect -4348 -1853 -4296 -1819
rect -4461 -1877 -4296 -1853
rect -4427 -1891 -4296 -1877
rect -4427 -1911 -4382 -1891
rect -4461 -1925 -4382 -1911
rect -4348 -1925 -4296 -1891
rect -4461 -1945 -4296 -1925
rect -4427 -1963 -4296 -1945
rect -4427 -1979 -4382 -1963
rect -4461 -1997 -4382 -1979
rect -4348 -1997 -4296 -1963
rect -4461 -2013 -4296 -1997
rect -4427 -2047 -4296 -2013
rect -4461 -2081 -4296 -2047
rect -4427 -2115 -4296 -2081
rect 2561 -687 2697 -653
rect 2561 -721 2731 -687
rect 2561 -755 2697 -721
rect 2561 -789 2731 -755
rect 2561 -823 2697 -789
rect 2561 -857 2731 -823
rect 2561 -891 2697 -857
rect 2561 -925 2731 -891
rect 2561 -959 2697 -925
rect 2561 -993 2731 -959
rect 2561 -1027 2697 -993
rect 2561 -1061 2731 -1027
rect 2561 -1095 2697 -1061
rect 2561 -1129 2731 -1095
rect 2561 -1163 2697 -1129
rect 2561 -1197 2731 -1163
rect 2561 -1231 2697 -1197
rect 2561 -1265 2731 -1231
rect 2561 -1299 2697 -1265
rect 2561 -1333 2731 -1299
rect 2561 -1367 2697 -1333
rect 2561 -1401 2731 -1367
rect 2561 -1435 2697 -1401
rect 2561 -1469 2731 -1435
rect 2561 -1503 2697 -1469
rect 2561 -1537 2731 -1503
rect 2561 -1571 2697 -1537
rect 2561 -1605 2731 -1571
rect 2561 -1639 2697 -1605
rect 2561 -1673 2731 -1639
rect 2561 -1707 2697 -1673
rect 2561 -1741 2731 -1707
rect 2561 -1775 2697 -1741
rect 2561 -1809 2731 -1775
rect 2561 -1843 2697 -1809
rect 2561 -1877 2731 -1843
rect 2561 -1911 2697 -1877
rect 2561 -1945 2731 -1911
rect 2561 -1979 2697 -1945
rect 2561 -2013 2731 -1979
rect 2561 -2047 2697 -2013
rect 2561 -2081 2731 -2047
rect -4461 -2149 -4296 -2115
rect -4427 -2183 -4296 -2149
rect -4461 -2217 -4296 -2183
rect -4427 -2251 -4296 -2217
rect -4461 -2285 -4296 -2251
rect -4427 -2319 -4296 -2285
rect -4461 -2353 -4296 -2319
rect -4427 -2387 -4296 -2353
rect -4461 -2421 -4296 -2387
rect -4427 -2455 -4296 -2421
rect -4461 -2489 -4296 -2455
rect -4427 -2523 -4296 -2489
rect -4461 -2557 -4296 -2523
rect -4427 -2591 -4296 -2557
rect -4461 -2618 -4296 -2591
rect -4461 -2625 -4375 -2618
rect -4427 -2652 -4375 -2625
rect -4341 -2652 -4296 -2618
rect -4427 -2659 -4296 -2652
rect -4461 -2690 -4296 -2659
rect -4461 -2693 -4375 -2690
rect -4427 -2724 -4375 -2693
rect -4341 -2724 -4296 -2690
rect -4427 -2727 -4296 -2724
rect -4461 -2761 -4296 -2727
rect -4427 -2762 -4296 -2761
rect -4427 -2795 -4375 -2762
rect -4461 -2796 -4375 -2795
rect -4341 -2796 -4296 -2762
rect -4461 -2829 -4296 -2796
rect -4427 -2834 -4296 -2829
rect -4427 -2863 -4375 -2834
rect -4461 -2868 -4375 -2863
rect -4341 -2868 -4296 -2834
rect -4461 -2897 -4296 -2868
rect -4427 -2906 -4296 -2897
rect -4427 -2931 -4375 -2906
rect -4461 -2940 -4375 -2931
rect -4341 -2940 -4296 -2906
rect -4461 -2965 -4296 -2940
rect -4427 -2978 -4296 -2965
rect -4427 -2999 -4375 -2978
rect -4461 -3012 -4375 -2999
rect -4341 -3012 -4296 -2978
rect -4461 -3033 -4296 -3012
rect -4427 -3050 -4296 -3033
rect -4427 -3067 -4375 -3050
rect -4461 -3084 -4375 -3067
rect -4341 -3084 -4296 -3050
rect -4461 -3101 -4296 -3084
rect -4427 -3122 -4296 -3101
rect -4427 -3135 -4375 -3122
rect -4461 -3156 -4375 -3135
rect -4341 -3156 -4296 -3122
rect -4461 -3169 -4296 -3156
rect -4427 -3194 -4296 -3169
rect -4427 -3203 -4375 -3194
rect -4461 -3228 -4375 -3203
rect -4341 -3228 -4296 -3194
rect -4461 -3237 -4296 -3228
rect -4427 -3266 -4296 -3237
rect -4427 -3271 -4375 -3266
rect -4461 -3300 -4375 -3271
rect -4341 -3300 -4296 -3266
rect -4461 -3305 -4296 -3300
rect -4427 -3338 -4296 -3305
rect -4427 -3339 -4375 -3338
rect -4461 -3372 -4375 -3339
rect -4341 -3372 -4296 -3338
rect -4461 -3373 -4296 -3372
rect -4427 -3407 -4296 -3373
rect -4461 -3410 -4296 -3407
rect -4461 -3441 -4375 -3410
rect -4427 -3444 -4375 -3441
rect -4341 -3444 -4296 -3410
rect -4427 -3475 -4296 -3444
rect -4461 -3482 -4296 -3475
rect -4461 -3509 -4375 -3482
rect -4427 -3516 -4375 -3509
rect -4341 -3516 -4296 -3482
rect -4427 -3543 -4296 -3516
rect -4461 -3554 -4296 -3543
rect -4461 -3577 -4375 -3554
rect -4427 -3588 -4375 -3577
rect -4341 -3588 -4296 -3554
rect -4427 -3611 -4296 -3588
rect -4175 -2108 -3937 -2103
rect -4175 -2167 2443 -2108
rect -4175 -2173 -3897 -2167
rect -4175 -2207 -4079 -2173
rect -4045 -2201 -3897 -2173
rect -3863 -2201 -3825 -2167
rect -3791 -2201 -3753 -2167
rect -3719 -2201 -3681 -2167
rect -3647 -2201 -3609 -2167
rect -3575 -2201 -3537 -2167
rect -3503 -2201 -3465 -2167
rect -3431 -2201 -3393 -2167
rect -3359 -2201 -3321 -2167
rect -3287 -2201 -3249 -2167
rect -3215 -2201 -3177 -2167
rect -3143 -2201 -3105 -2167
rect -3071 -2201 -3033 -2167
rect -2999 -2201 -2961 -2167
rect -2927 -2201 -2889 -2167
rect -2855 -2201 -2817 -2167
rect -2783 -2201 -2745 -2167
rect -2711 -2201 -2673 -2167
rect -2639 -2201 -2601 -2167
rect -2567 -2201 -2529 -2167
rect -2495 -2201 -2457 -2167
rect -2423 -2201 -2385 -2167
rect -2351 -2201 -2313 -2167
rect -2279 -2201 -2241 -2167
rect -2207 -2201 -2169 -2167
rect -2135 -2201 -2097 -2167
rect -2063 -2201 -2025 -2167
rect -1991 -2201 -1953 -2167
rect -1919 -2201 -1881 -2167
rect -1847 -2201 -1809 -2167
rect -1775 -2201 -1737 -2167
rect -1703 -2201 -1665 -2167
rect -1631 -2201 -1593 -2167
rect -1559 -2201 -1521 -2167
rect -1487 -2201 -1449 -2167
rect -1415 -2201 -1377 -2167
rect -1343 -2201 -1305 -2167
rect -1271 -2201 -1233 -2167
rect -1199 -2201 -1161 -2167
rect -1127 -2201 -1089 -2167
rect -1055 -2201 -1017 -2167
rect -983 -2201 -945 -2167
rect -911 -2201 -873 -2167
rect -839 -2201 -801 -2167
rect -767 -2201 -729 -2167
rect -695 -2201 -657 -2167
rect -623 -2201 -585 -2167
rect -551 -2201 -513 -2167
rect -479 -2201 -441 -2167
rect -407 -2201 -369 -2167
rect -335 -2201 -297 -2167
rect -263 -2201 -225 -2167
rect -191 -2201 -153 -2167
rect -119 -2201 -81 -2167
rect -47 -2201 -9 -2167
rect 25 -2201 63 -2167
rect 97 -2201 135 -2167
rect 169 -2201 207 -2167
rect 241 -2201 279 -2167
rect 313 -2201 351 -2167
rect 385 -2201 423 -2167
rect 457 -2201 495 -2167
rect 529 -2201 567 -2167
rect 601 -2201 639 -2167
rect 673 -2201 711 -2167
rect 745 -2201 783 -2167
rect 817 -2201 855 -2167
rect 889 -2201 927 -2167
rect 961 -2201 999 -2167
rect 1033 -2201 1071 -2167
rect 1105 -2201 1143 -2167
rect 1177 -2201 1215 -2167
rect 1249 -2201 1287 -2167
rect 1321 -2201 1359 -2167
rect 1393 -2201 1431 -2167
rect 1465 -2201 1503 -2167
rect 1537 -2201 1575 -2167
rect 1609 -2201 1647 -2167
rect 1681 -2201 1719 -2167
rect 1753 -2201 1791 -2167
rect 1825 -2201 1863 -2167
rect 1897 -2201 1935 -2167
rect 1969 -2201 2007 -2167
rect 2041 -2201 2079 -2167
rect 2113 -2201 2151 -2167
rect 2185 -2201 2223 -2167
rect 2257 -2201 2295 -2167
rect 2329 -2201 2443 -2167
rect -4045 -2207 2443 -2201
rect -4175 -2245 2443 -2207
rect -4175 -2279 -4079 -2245
rect -4045 -2259 2443 -2245
rect -4045 -2279 -3937 -2259
rect -4175 -2317 -3937 -2279
rect -4175 -2351 -4079 -2317
rect -4045 -2351 -3937 -2317
rect -4175 -2389 -3937 -2351
rect -4175 -2423 -4079 -2389
rect -4045 -2423 -3937 -2389
rect -4175 -2461 -3937 -2423
rect -4175 -2495 -4079 -2461
rect -4045 -2495 -3937 -2461
rect -4175 -2533 -3937 -2495
rect -4175 -2567 -4079 -2533
rect -4045 -2567 -3937 -2533
rect -4175 -2605 -3937 -2567
rect -4175 -2639 -4079 -2605
rect -4045 -2639 -3937 -2605
rect -4175 -2677 -3937 -2639
rect -4175 -2711 -4079 -2677
rect -4045 -2711 -3937 -2677
rect -4175 -2749 -3937 -2711
rect -4175 -2783 -4079 -2749
rect -4045 -2783 -3937 -2749
rect -4175 -2821 -3937 -2783
rect -4175 -2855 -4079 -2821
rect -4045 -2855 -3937 -2821
rect -4175 -2893 -3937 -2855
rect -4175 -2927 -4079 -2893
rect -4045 -2927 -3937 -2893
rect -4175 -2965 -3937 -2927
rect -4175 -2999 -4079 -2965
rect -4045 -2999 -3937 -2965
rect -4175 -3037 -3937 -2999
rect -4175 -3071 -4079 -3037
rect -4045 -3071 -3937 -3037
rect -4175 -3109 -3937 -3071
rect -4175 -3143 -4079 -3109
rect -4045 -3143 -3937 -3109
rect -4175 -3181 -3937 -3143
rect -4175 -3215 -4079 -3181
rect -4045 -3215 -3937 -3181
rect -4175 -3253 -3937 -3215
rect -4175 -3287 -4079 -3253
rect -4045 -3287 -3937 -3253
rect -4175 -3325 -3937 -3287
rect -4175 -3359 -4079 -3325
rect -4045 -3359 -3937 -3325
rect -4175 -3397 -3937 -3359
rect -4175 -3431 -4079 -3397
rect -4045 -3431 -3937 -3397
rect -4175 -3469 -3937 -3431
rect -4175 -3503 -4079 -3469
rect -4045 -3503 -3937 -3469
rect -4175 -3508 -3937 -3503
rect 2153 -2503 2443 -2259
rect 2153 -2537 2327 -2503
rect 2361 -2537 2443 -2503
rect 2153 -2575 2443 -2537
rect 2153 -2609 2327 -2575
rect 2361 -2609 2443 -2575
rect 2153 -2647 2443 -2609
rect 2153 -2681 2327 -2647
rect 2361 -2681 2443 -2647
rect 2153 -2719 2443 -2681
rect 2153 -2753 2327 -2719
rect 2361 -2753 2443 -2719
rect 2153 -2791 2443 -2753
rect 2153 -2825 2327 -2791
rect 2361 -2825 2443 -2791
rect 2153 -2863 2443 -2825
rect 2153 -2897 2327 -2863
rect 2361 -2897 2443 -2863
rect 2153 -2935 2443 -2897
rect 2153 -2969 2327 -2935
rect 2361 -2969 2443 -2935
rect 2153 -3007 2443 -2969
rect 2153 -3041 2327 -3007
rect 2361 -3041 2443 -3007
rect 2153 -3079 2443 -3041
rect 2153 -3113 2327 -3079
rect 2361 -3113 2443 -3079
rect 2153 -3151 2443 -3113
rect 2153 -3185 2327 -3151
rect 2361 -3185 2443 -3151
rect 2153 -3223 2443 -3185
rect 2153 -3257 2327 -3223
rect 2361 -3257 2443 -3223
rect 2153 -3295 2443 -3257
rect 2153 -3329 2327 -3295
rect 2361 -3329 2443 -3295
rect 2153 -3367 2443 -3329
rect 2153 -3401 2327 -3367
rect 2361 -3401 2443 -3367
rect 2153 -3439 2443 -3401
rect 2153 -3473 2327 -3439
rect 2361 -3473 2443 -3439
rect 2153 -3508 2443 -3473
rect -4175 -3511 2443 -3508
rect -4175 -3545 2327 -3511
rect 2361 -3545 2443 -3511
rect -4175 -3548 2443 -3545
rect -4175 -3582 -3970 -3548
rect -3936 -3582 -3898 -3548
rect -3864 -3582 -3826 -3548
rect -3792 -3582 -3754 -3548
rect -3720 -3582 -3682 -3548
rect -3648 -3582 -3610 -3548
rect -3576 -3582 -3538 -3548
rect -3504 -3582 -3466 -3548
rect -3432 -3582 -3394 -3548
rect -3360 -3582 -3322 -3548
rect -3288 -3582 -3250 -3548
rect -3216 -3582 -3178 -3548
rect -3144 -3582 -3106 -3548
rect -3072 -3582 -3034 -3548
rect -3000 -3582 -2962 -3548
rect -2928 -3582 -2890 -3548
rect -2856 -3582 -2818 -3548
rect -2784 -3582 -2746 -3548
rect -2712 -3582 -2674 -3548
rect -2640 -3582 -2602 -3548
rect -2568 -3582 -2530 -3548
rect -2496 -3582 -2458 -3548
rect -2424 -3582 -2386 -3548
rect -2352 -3582 -2314 -3548
rect -2280 -3582 -2242 -3548
rect -2208 -3582 -2170 -3548
rect -2136 -3582 -2098 -3548
rect -2064 -3582 -2026 -3548
rect -1992 -3582 -1954 -3548
rect -1920 -3582 -1882 -3548
rect -1848 -3582 -1810 -3548
rect -1776 -3582 -1738 -3548
rect -1704 -3582 -1666 -3548
rect -1632 -3582 -1594 -3548
rect -1560 -3582 -1522 -3548
rect -1488 -3582 -1450 -3548
rect -1416 -3582 -1378 -3548
rect -1344 -3582 -1306 -3548
rect -1272 -3582 -1234 -3548
rect -1200 -3582 -1162 -3548
rect -1128 -3582 -1090 -3548
rect -1056 -3582 -1018 -3548
rect -984 -3582 -946 -3548
rect -912 -3582 -874 -3548
rect -840 -3582 -802 -3548
rect -768 -3582 -730 -3548
rect -696 -3582 -658 -3548
rect -624 -3582 -586 -3548
rect -552 -3582 -514 -3548
rect -480 -3582 -442 -3548
rect -408 -3582 -370 -3548
rect -336 -3582 -298 -3548
rect -264 -3582 -226 -3548
rect -192 -3582 -154 -3548
rect -120 -3582 -82 -3548
rect -48 -3582 -10 -3548
rect 24 -3582 62 -3548
rect 96 -3582 134 -3548
rect 168 -3582 206 -3548
rect 240 -3582 278 -3548
rect 312 -3582 350 -3548
rect 384 -3582 422 -3548
rect 456 -3582 494 -3548
rect 528 -3582 566 -3548
rect 600 -3582 638 -3548
rect 672 -3582 710 -3548
rect 744 -3582 782 -3548
rect 816 -3582 854 -3548
rect 888 -3582 926 -3548
rect 960 -3582 998 -3548
rect 1032 -3582 1070 -3548
rect 1104 -3582 1142 -3548
rect 1176 -3582 1214 -3548
rect 1248 -3582 1286 -3548
rect 1320 -3582 1358 -3548
rect 1392 -3582 1430 -3548
rect 1464 -3582 1502 -3548
rect 1536 -3582 1574 -3548
rect 1608 -3582 1646 -3548
rect 1680 -3582 1718 -3548
rect 1752 -3582 1790 -3548
rect 1824 -3582 1862 -3548
rect 1896 -3582 1934 -3548
rect 1968 -3582 2006 -3548
rect 2040 -3582 2078 -3548
rect 2112 -3582 2150 -3548
rect 2184 -3582 2222 -3548
rect 2256 -3582 2443 -3548
rect -4175 -3606 2443 -3582
rect 2561 -2115 2697 -2081
rect 2561 -2149 2731 -2115
rect 2561 -2183 2697 -2149
rect 2561 -2217 2731 -2183
rect 2561 -2251 2697 -2217
rect 2561 -2285 2731 -2251
rect 2561 -2319 2697 -2285
rect 2561 -2353 2731 -2319
rect 2561 -2387 2697 -2353
rect 2561 -2421 2731 -2387
rect 2561 -2455 2697 -2421
rect 2561 -2489 2731 -2455
rect 2561 -2500 2697 -2489
rect 2561 -2534 2610 -2500
rect 2644 -2523 2697 -2500
rect 2644 -2534 2731 -2523
rect 2561 -2557 2731 -2534
rect 2561 -2572 2697 -2557
rect 2561 -2606 2610 -2572
rect 2644 -2591 2697 -2572
rect 2644 -2606 2731 -2591
rect 2561 -2625 2731 -2606
rect 2561 -2644 2697 -2625
rect 2561 -2678 2610 -2644
rect 2644 -2659 2697 -2644
rect 2644 -2678 2731 -2659
rect 2561 -2693 2731 -2678
rect 2561 -2716 2697 -2693
rect 2561 -2750 2610 -2716
rect 2644 -2727 2697 -2716
rect 2644 -2750 2731 -2727
rect 2561 -2761 2731 -2750
rect 2561 -2788 2697 -2761
rect 2561 -2822 2610 -2788
rect 2644 -2795 2697 -2788
rect 2644 -2822 2731 -2795
rect 2561 -2829 2731 -2822
rect 2561 -2860 2697 -2829
rect 2561 -2894 2610 -2860
rect 2644 -2863 2697 -2860
rect 2644 -2894 2731 -2863
rect 2561 -2897 2731 -2894
rect 2561 -2931 2697 -2897
rect 2561 -2932 2731 -2931
rect 2561 -2966 2610 -2932
rect 2644 -2965 2731 -2932
rect 2644 -2966 2697 -2965
rect 2561 -2999 2697 -2966
rect 2561 -3004 2731 -2999
rect 2561 -3038 2610 -3004
rect 2644 -3033 2731 -3004
rect 2644 -3038 2697 -3033
rect 2561 -3067 2697 -3038
rect 2561 -3076 2731 -3067
rect 2561 -3110 2610 -3076
rect 2644 -3101 2731 -3076
rect 2644 -3110 2697 -3101
rect 2561 -3135 2697 -3110
rect 2561 -3148 2731 -3135
rect 2561 -3182 2610 -3148
rect 2644 -3169 2731 -3148
rect 2644 -3182 2697 -3169
rect 2561 -3203 2697 -3182
rect 2561 -3231 2731 -3203
rect 2561 -3481 2576 -3231
rect 2682 -3237 2731 -3231
rect 2682 -3271 2697 -3237
rect 2682 -3305 2731 -3271
rect 2682 -3339 2697 -3305
rect 2682 -3373 2731 -3339
rect 2682 -3407 2697 -3373
rect 2682 -3441 2731 -3407
rect 2682 -3475 2697 -3441
rect 2682 -3481 2731 -3475
rect 2561 -3509 2731 -3481
rect 2561 -3543 2697 -3509
rect 2561 -3577 2731 -3543
rect -4461 -3645 -4296 -3611
rect -4427 -3654 -4296 -3645
rect 2561 -3611 2697 -3577
rect 2561 -3645 2731 -3611
rect 2561 -3654 2697 -3645
rect -4427 -3679 2697 -3654
rect -4461 -3696 2731 -3679
rect -4461 -3713 -4371 -3696
rect -4427 -3730 -4371 -3713
rect -4337 -3730 -4299 -3696
rect -4265 -3730 -4227 -3696
rect -4193 -3730 -4155 -3696
rect -4121 -3730 -4083 -3696
rect -4049 -3730 -4011 -3696
rect -3977 -3730 -3939 -3696
rect -3905 -3730 -3867 -3696
rect -3833 -3730 -3795 -3696
rect -3761 -3730 -3723 -3696
rect -3689 -3730 -3651 -3696
rect -3617 -3730 -3579 -3696
rect -3545 -3730 -3507 -3696
rect -3473 -3730 -3435 -3696
rect -3401 -3730 -3363 -3696
rect -3329 -3730 -3291 -3696
rect -3257 -3730 -3219 -3696
rect -3185 -3730 -3147 -3696
rect -3113 -3730 -3075 -3696
rect -3041 -3730 -3003 -3696
rect -2969 -3730 -2931 -3696
rect -2897 -3730 -2859 -3696
rect -2825 -3730 -2787 -3696
rect -2753 -3730 -2715 -3696
rect -2681 -3730 -2643 -3696
rect -2609 -3730 -2571 -3696
rect -2537 -3730 -2499 -3696
rect -2465 -3730 -2427 -3696
rect -2393 -3730 -2355 -3696
rect -2321 -3730 -2283 -3696
rect -2249 -3730 -2211 -3696
rect -2177 -3730 -2139 -3696
rect -2105 -3730 -2067 -3696
rect -2033 -3730 -1995 -3696
rect -1961 -3730 -1923 -3696
rect -1889 -3730 -1851 -3696
rect -1817 -3730 -1779 -3696
rect -1745 -3730 -1707 -3696
rect -1673 -3730 -1635 -3696
rect -1601 -3730 -1563 -3696
rect -1529 -3730 -1491 -3696
rect -1457 -3730 -1419 -3696
rect -1385 -3730 -1347 -3696
rect -1313 -3730 -1275 -3696
rect -1241 -3730 -1203 -3696
rect -1169 -3730 -1131 -3696
rect -1097 -3730 -1059 -3696
rect -1025 -3730 -987 -3696
rect -953 -3730 -915 -3696
rect -881 -3730 -843 -3696
rect -809 -3730 -771 -3696
rect -737 -3730 -699 -3696
rect -665 -3730 -627 -3696
rect -593 -3730 -555 -3696
rect -521 -3730 -483 -3696
rect -449 -3730 -411 -3696
rect -377 -3730 -339 -3696
rect -305 -3730 -267 -3696
rect -233 -3730 -195 -3696
rect -161 -3730 -123 -3696
rect -89 -3730 -51 -3696
rect -17 -3730 21 -3696
rect 55 -3730 93 -3696
rect 127 -3730 165 -3696
rect 199 -3730 237 -3696
rect 271 -3730 309 -3696
rect 343 -3730 381 -3696
rect 415 -3730 453 -3696
rect 487 -3730 525 -3696
rect 559 -3730 597 -3696
rect 631 -3730 669 -3696
rect 703 -3730 741 -3696
rect 775 -3730 813 -3696
rect 847 -3730 885 -3696
rect 919 -3730 957 -3696
rect 991 -3730 1029 -3696
rect 1063 -3730 1101 -3696
rect 1135 -3730 1173 -3696
rect 1207 -3730 1245 -3696
rect 1279 -3730 1317 -3696
rect 1351 -3730 1389 -3696
rect 1423 -3730 1461 -3696
rect 1495 -3730 1533 -3696
rect 1567 -3730 1605 -3696
rect 1639 -3730 1677 -3696
rect 1711 -3730 1749 -3696
rect 1783 -3730 1821 -3696
rect 1855 -3730 1893 -3696
rect 1927 -3730 1965 -3696
rect 1999 -3730 2037 -3696
rect 2071 -3730 2109 -3696
rect 2143 -3730 2181 -3696
rect 2215 -3730 2253 -3696
rect 2287 -3730 2325 -3696
rect 2359 -3730 2397 -3696
rect 2431 -3730 2469 -3696
rect 2503 -3730 2541 -3696
rect 2575 -3730 2613 -3696
rect 2647 -3713 2731 -3696
rect 2647 -3730 2697 -3713
rect -4427 -3747 2697 -3730
rect -4461 -3781 2731 -3747
rect -4461 -3815 -4384 -3781
rect -4350 -3815 -4316 -3781
rect -4282 -3815 -4248 -3781
rect -4214 -3815 -4180 -3781
rect -4146 -3815 -4112 -3781
rect -4078 -3815 -4044 -3781
rect -4010 -3815 -3976 -3781
rect -3942 -3815 -3908 -3781
rect -3874 -3815 -3840 -3781
rect -3806 -3815 -3772 -3781
rect -3738 -3815 -3704 -3781
rect -3670 -3815 -3636 -3781
rect -3602 -3815 -3568 -3781
rect -3534 -3815 -3500 -3781
rect -3466 -3815 -3432 -3781
rect -3398 -3815 -3364 -3781
rect -3330 -3815 -3296 -3781
rect -3262 -3815 -3228 -3781
rect -3194 -3815 -3160 -3781
rect -3126 -3815 -3092 -3781
rect -3058 -3815 -3024 -3781
rect -2990 -3815 -2956 -3781
rect -2922 -3815 -2888 -3781
rect -2854 -3815 -2820 -3781
rect -2786 -3815 -2752 -3781
rect -2718 -3815 -2684 -3781
rect -2650 -3815 -2616 -3781
rect -2582 -3815 -2548 -3781
rect -2514 -3815 -2480 -3781
rect -2446 -3815 -2412 -3781
rect -2378 -3815 -2344 -3781
rect -2310 -3815 -2276 -3781
rect -2242 -3815 -2208 -3781
rect -2174 -3815 -2140 -3781
rect -2106 -3815 -2072 -3781
rect -2038 -3815 -2004 -3781
rect -1970 -3815 -1936 -3781
rect -1902 -3815 -1868 -3781
rect -1834 -3815 -1800 -3781
rect -1766 -3815 -1732 -3781
rect -1698 -3815 -1664 -3781
rect -1630 -3815 -1596 -3781
rect -1562 -3815 -1528 -3781
rect -1494 -3815 -1460 -3781
rect -1426 -3815 -1392 -3781
rect -1358 -3815 -1324 -3781
rect -1290 -3815 -1256 -3781
rect -1222 -3815 -1188 -3781
rect -1154 -3815 -1120 -3781
rect -1086 -3815 -1052 -3781
rect -1018 -3815 -984 -3781
rect -950 -3815 -916 -3781
rect -882 -3815 -848 -3781
rect -814 -3815 -780 -3781
rect -746 -3815 -712 -3781
rect -678 -3815 -644 -3781
rect -610 -3815 -576 -3781
rect -542 -3815 -508 -3781
rect -474 -3815 -440 -3781
rect -406 -3815 -372 -3781
rect -338 -3815 -304 -3781
rect -270 -3815 -236 -3781
rect -202 -3815 -168 -3781
rect -134 -3815 -100 -3781
rect -66 -3815 -32 -3781
rect 2 -3815 36 -3781
rect 70 -3815 104 -3781
rect 138 -3815 172 -3781
rect 206 -3815 240 -3781
rect 274 -3815 308 -3781
rect 342 -3815 376 -3781
rect 410 -3815 444 -3781
rect 478 -3815 512 -3781
rect 546 -3815 580 -3781
rect 614 -3815 648 -3781
rect 682 -3815 716 -3781
rect 750 -3815 784 -3781
rect 818 -3815 852 -3781
rect 886 -3815 920 -3781
rect 954 -3815 988 -3781
rect 1022 -3815 1056 -3781
rect 1090 -3815 1124 -3781
rect 1158 -3815 1192 -3781
rect 1226 -3815 1260 -3781
rect 1294 -3815 1328 -3781
rect 1362 -3815 1396 -3781
rect 1430 -3815 1464 -3781
rect 1498 -3815 1532 -3781
rect 1566 -3815 1600 -3781
rect 1634 -3815 1668 -3781
rect 1702 -3815 1736 -3781
rect 1770 -3815 1804 -3781
rect 1838 -3815 1872 -3781
rect 1906 -3815 1940 -3781
rect 1974 -3815 2008 -3781
rect 2042 -3815 2076 -3781
rect 2110 -3815 2144 -3781
rect 2178 -3815 2212 -3781
rect 2246 -3815 2280 -3781
rect 2314 -3815 2348 -3781
rect 2382 -3815 2416 -3781
rect 2450 -3815 2484 -3781
rect 2518 -3815 2552 -3781
rect 2586 -3815 2620 -3781
rect 2654 -3815 2731 -3781
<< viali >>
rect -4317 6364 2629 6470
rect -4318 6262 -4284 6296
rect -4318 6190 -4284 6224
rect -4318 6118 -4284 6152
rect -4318 6046 -4284 6080
rect -4318 5974 -4284 6008
rect -4318 5902 -4284 5936
rect -4318 5830 -4284 5864
rect -4318 5758 -4284 5792
rect -4318 5686 -4284 5720
rect -4318 5614 -4284 5648
rect -4318 5542 -4284 5576
rect -4318 5470 -4284 5504
rect -4318 5398 -4284 5432
rect -4318 5326 -4284 5360
rect -4318 5254 -4284 5288
rect -4318 5182 -4284 5216
rect -4318 5110 -4284 5144
rect -4318 5038 -4284 5072
rect -4318 4966 -4284 5000
rect -4318 4894 -4284 4928
rect -4318 4822 -4284 4856
rect -4318 4750 -4284 4784
rect -4318 4678 -4284 4712
rect -4318 4606 -4284 4640
rect -4318 4534 -4284 4568
rect -4318 4462 -4284 4496
rect -4318 4390 -4284 4424
rect -4318 4318 -4284 4352
rect -4318 4246 -4284 4280
rect -4318 4174 -4284 4208
rect -4148 3892 -4114 3926
rect -4076 3892 -4042 3926
rect -4004 3892 -3970 3926
rect -3932 3892 -3898 3926
rect -3860 3892 -3826 3926
rect -3788 3892 -3754 3926
rect -3716 3892 -3682 3926
rect -3644 3892 -3610 3926
rect -3572 3892 -3538 3926
rect -3500 3892 -3466 3926
rect -3428 3892 -3394 3926
rect -3356 3892 -3322 3926
rect -3284 3892 -3250 3926
rect -3212 3892 -3178 3926
rect -3140 3892 -3106 3926
rect -3068 3892 -3034 3926
rect -2996 3892 -2962 3926
rect -2924 3892 -2890 3926
rect -2852 3892 -2818 3926
rect -2780 3892 -2746 3926
rect -2708 3892 -2674 3926
rect -2636 3892 -2602 3926
rect -2564 3892 -2530 3926
rect -2492 3892 -2458 3926
rect -2420 3892 -2386 3926
rect -2348 3892 -2314 3926
rect -2276 3892 -2242 3926
rect -2204 3892 -2170 3926
rect -2132 3892 -2098 3926
rect -2060 3892 -2026 3926
rect -1988 3892 -1954 3926
rect -1916 3892 -1882 3926
rect -1844 3892 -1810 3926
rect -1772 3892 -1738 3926
rect -1700 3892 -1666 3926
rect -1628 3892 -1594 3926
rect -1556 3892 -1522 3926
rect -1484 3892 -1450 3926
rect -1412 3892 -1378 3926
rect -1340 3892 -1306 3926
rect -1268 3892 -1234 3926
rect -1196 3892 -1162 3926
rect -1124 3892 -1090 3926
rect -1052 3892 -1018 3926
rect -980 3892 -946 3926
rect -908 3892 -874 3926
rect -836 3892 -802 3926
rect -764 3892 -730 3926
rect -692 3892 -658 3926
rect -620 3892 -586 3926
rect -548 3892 -514 3926
rect -476 3892 -442 3926
rect -404 3892 -370 3926
rect -332 3892 -298 3926
rect -260 3892 -226 3926
rect -188 3892 -154 3926
rect -116 3892 -82 3926
rect -44 3892 -10 3926
rect 28 3892 62 3926
rect 100 3892 134 3926
rect 172 3892 206 3926
rect 244 3892 278 3926
rect 316 3892 350 3926
rect 388 3892 422 3926
rect 460 3892 494 3926
rect 532 3892 566 3926
rect 604 3892 638 3926
rect 676 3892 710 3926
rect 748 3892 782 3926
rect 820 3892 854 3926
rect 892 3892 926 3926
rect 964 3892 998 3926
rect 1036 3892 1070 3926
rect 1108 3892 1142 3926
rect 1180 3892 1214 3926
rect 1252 3892 1286 3926
rect 1324 3892 1358 3926
rect 1396 3892 1430 3926
rect 1468 3892 1502 3926
rect 1540 3892 1574 3926
rect 1612 3892 1646 3926
rect 1684 3892 1718 3926
rect 1756 3892 1790 3926
rect 1828 3892 1862 3926
rect 1900 3892 1934 3926
rect 1972 3892 2006 3926
rect 2044 3892 2078 3926
rect 2116 3892 2150 3926
rect 2188 3892 2222 3926
rect 2260 3892 2294 3926
rect 2332 3892 2366 3926
rect 2404 3892 2438 3926
rect -4035 1221 -3857 1399
rect -4342 929 -4164 1179
rect -3397 555 -3291 1381
rect -3193 1260 1305 1366
rect 1404 502 1510 1400
rect 2148 1223 2326 1401
rect -4382 -701 -4348 -667
rect -4105 -523 -3999 15
rect -3509 -451 -3403 15
rect -3652 -617 -3618 -583
rect -3580 -617 -3546 -583
rect -3508 -617 -3474 -583
rect -3436 -617 -3402 -583
rect -3364 -617 -3330 -583
rect -3292 -617 -3258 -583
rect -3220 -617 -3186 -583
rect -3148 -617 -3114 -583
rect -3076 -617 -3042 -583
rect -3004 -617 -2970 -583
rect -2932 -617 -2898 -583
rect -2860 -617 -2826 -583
rect -2788 -617 -2754 -583
rect -2716 -617 -2682 -583
rect -2644 -617 -2610 -583
rect -2572 -617 -2538 -583
rect -2500 -617 -2466 -583
rect -2428 -617 -2394 -583
rect -2356 -617 -2322 -583
rect -2284 -617 -2250 -583
rect -2212 -617 -2178 -583
rect -2140 -617 -2106 -583
rect -2068 -617 -2034 -583
rect -1996 -617 -1962 -583
rect -1924 -617 -1890 -583
rect -1852 -617 -1818 -583
rect -1780 -617 -1746 -583
rect -1708 -617 -1674 -583
rect -1636 -617 -1602 -583
rect -1564 -617 -1530 -583
rect -1492 -617 -1458 -583
rect -1420 -617 -1386 -583
rect -1348 -617 -1314 -583
rect -1276 -617 -1242 -583
rect -1204 -617 -1170 -583
rect -1132 -617 -1098 -583
rect -1060 -617 -1026 -583
rect -988 -617 -954 -583
rect -916 -617 -882 -583
rect -844 -617 -810 -583
rect -772 -617 -738 -583
rect -700 -617 -666 -583
rect -628 -617 -594 -583
rect -556 -617 -522 -583
rect -484 -617 -450 -583
rect -412 -617 -378 -583
rect -340 -617 -306 -583
rect -268 -617 -234 -583
rect -196 -617 -162 -583
rect -124 -617 -90 -583
rect -52 -617 -18 -583
rect 20 -617 54 -583
rect 92 -617 126 -583
rect 164 -617 198 -583
rect 236 -617 270 -583
rect 308 -617 342 -583
rect 380 -617 414 -583
rect 452 -617 486 -583
rect 524 -617 558 -583
rect 596 -617 630 -583
rect 668 -617 702 -583
rect 740 -617 774 -583
rect 812 -617 846 -583
rect 884 -617 918 -583
rect 956 -617 990 -583
rect 1028 -617 1062 -583
rect 1100 -617 1134 -583
rect 1172 -617 1206 -583
rect 1244 -617 1278 -583
rect 1316 -617 1350 -583
rect 1388 -617 1422 -583
rect 1460 -617 1494 -583
rect 1532 -617 1566 -583
rect 1604 -617 1638 -583
rect 1676 -617 1710 -583
rect 1748 -617 1782 -583
rect 1820 -617 1854 -583
rect 1892 -617 1926 -583
rect 1964 -617 1998 -583
rect 2036 -617 2070 -583
rect 2108 -617 2142 -583
rect 2180 -617 2214 -583
rect -4382 -773 -4348 -739
rect -4382 -845 -4348 -811
rect -4382 -917 -4348 -883
rect -4382 -989 -4348 -955
rect -4382 -1061 -4348 -1027
rect -4382 -1133 -4348 -1099
rect -4382 -1205 -4348 -1171
rect -4382 -1277 -4348 -1243
rect -4382 -1349 -4348 -1315
rect -4382 -1421 -4348 -1387
rect -4382 -1493 -4348 -1459
rect -4382 -1565 -4348 -1531
rect -4382 -1637 -4348 -1603
rect -4382 -1709 -4348 -1675
rect -4382 -1781 -4348 -1747
rect -4382 -1853 -4348 -1819
rect -4382 -1925 -4348 -1891
rect -4382 -1997 -4348 -1963
rect -4375 -2652 -4341 -2618
rect -4375 -2724 -4341 -2690
rect -4375 -2796 -4341 -2762
rect -4375 -2868 -4341 -2834
rect -4375 -2940 -4341 -2906
rect -4375 -3012 -4341 -2978
rect -4375 -3084 -4341 -3050
rect -4375 -3156 -4341 -3122
rect -4375 -3228 -4341 -3194
rect -4375 -3300 -4341 -3266
rect -4375 -3372 -4341 -3338
rect -4375 -3444 -4341 -3410
rect -4375 -3516 -4341 -3482
rect -4375 -3588 -4341 -3554
rect -4079 -2207 -4045 -2173
rect -3897 -2201 -3863 -2167
rect -3825 -2201 -3791 -2167
rect -3753 -2201 -3719 -2167
rect -3681 -2201 -3647 -2167
rect -3609 -2201 -3575 -2167
rect -3537 -2201 -3503 -2167
rect -3465 -2201 -3431 -2167
rect -3393 -2201 -3359 -2167
rect -3321 -2201 -3287 -2167
rect -3249 -2201 -3215 -2167
rect -3177 -2201 -3143 -2167
rect -3105 -2201 -3071 -2167
rect -3033 -2201 -2999 -2167
rect -2961 -2201 -2927 -2167
rect -2889 -2201 -2855 -2167
rect -2817 -2201 -2783 -2167
rect -2745 -2201 -2711 -2167
rect -2673 -2201 -2639 -2167
rect -2601 -2201 -2567 -2167
rect -2529 -2201 -2495 -2167
rect -2457 -2201 -2423 -2167
rect -2385 -2201 -2351 -2167
rect -2313 -2201 -2279 -2167
rect -2241 -2201 -2207 -2167
rect -2169 -2201 -2135 -2167
rect -2097 -2201 -2063 -2167
rect -2025 -2201 -1991 -2167
rect -1953 -2201 -1919 -2167
rect -1881 -2201 -1847 -2167
rect -1809 -2201 -1775 -2167
rect -1737 -2201 -1703 -2167
rect -1665 -2201 -1631 -2167
rect -1593 -2201 -1559 -2167
rect -1521 -2201 -1487 -2167
rect -1449 -2201 -1415 -2167
rect -1377 -2201 -1343 -2167
rect -1305 -2201 -1271 -2167
rect -1233 -2201 -1199 -2167
rect -1161 -2201 -1127 -2167
rect -1089 -2201 -1055 -2167
rect -1017 -2201 -983 -2167
rect -945 -2201 -911 -2167
rect -873 -2201 -839 -2167
rect -801 -2201 -767 -2167
rect -729 -2201 -695 -2167
rect -657 -2201 -623 -2167
rect -585 -2201 -551 -2167
rect -513 -2201 -479 -2167
rect -441 -2201 -407 -2167
rect -369 -2201 -335 -2167
rect -297 -2201 -263 -2167
rect -225 -2201 -191 -2167
rect -153 -2201 -119 -2167
rect -81 -2201 -47 -2167
rect -9 -2201 25 -2167
rect 63 -2201 97 -2167
rect 135 -2201 169 -2167
rect 207 -2201 241 -2167
rect 279 -2201 313 -2167
rect 351 -2201 385 -2167
rect 423 -2201 457 -2167
rect 495 -2201 529 -2167
rect 567 -2201 601 -2167
rect 639 -2201 673 -2167
rect 711 -2201 745 -2167
rect 783 -2201 817 -2167
rect 855 -2201 889 -2167
rect 927 -2201 961 -2167
rect 999 -2201 1033 -2167
rect 1071 -2201 1105 -2167
rect 1143 -2201 1177 -2167
rect 1215 -2201 1249 -2167
rect 1287 -2201 1321 -2167
rect 1359 -2201 1393 -2167
rect 1431 -2201 1465 -2167
rect 1503 -2201 1537 -2167
rect 1575 -2201 1609 -2167
rect 1647 -2201 1681 -2167
rect 1719 -2201 1753 -2167
rect 1791 -2201 1825 -2167
rect 1863 -2201 1897 -2167
rect 1935 -2201 1969 -2167
rect 2007 -2201 2041 -2167
rect 2079 -2201 2113 -2167
rect 2151 -2201 2185 -2167
rect 2223 -2201 2257 -2167
rect 2295 -2201 2329 -2167
rect -4079 -2279 -4045 -2245
rect -4079 -2351 -4045 -2317
rect -4079 -2423 -4045 -2389
rect -4079 -2495 -4045 -2461
rect -4079 -2567 -4045 -2533
rect -4079 -2639 -4045 -2605
rect -4079 -2711 -4045 -2677
rect -4079 -2783 -4045 -2749
rect -4079 -2855 -4045 -2821
rect -4079 -2927 -4045 -2893
rect -4079 -2999 -4045 -2965
rect -4079 -3071 -4045 -3037
rect -4079 -3143 -4045 -3109
rect -4079 -3215 -4045 -3181
rect -4079 -3287 -4045 -3253
rect -4079 -3359 -4045 -3325
rect -4079 -3431 -4045 -3397
rect -4079 -3503 -4045 -3469
rect 2327 -2537 2361 -2503
rect 2327 -2609 2361 -2575
rect 2327 -2681 2361 -2647
rect 2327 -2753 2361 -2719
rect 2327 -2825 2361 -2791
rect 2327 -2897 2361 -2863
rect 2327 -2969 2361 -2935
rect 2327 -3041 2361 -3007
rect 2327 -3113 2361 -3079
rect 2327 -3185 2361 -3151
rect 2327 -3257 2361 -3223
rect 2327 -3329 2361 -3295
rect 2327 -3401 2361 -3367
rect 2327 -3473 2361 -3439
rect 2327 -3545 2361 -3511
rect -3970 -3582 -3936 -3548
rect -3898 -3582 -3864 -3548
rect -3826 -3582 -3792 -3548
rect -3754 -3582 -3720 -3548
rect -3682 -3582 -3648 -3548
rect -3610 -3582 -3576 -3548
rect -3538 -3582 -3504 -3548
rect -3466 -3582 -3432 -3548
rect -3394 -3582 -3360 -3548
rect -3322 -3582 -3288 -3548
rect -3250 -3582 -3216 -3548
rect -3178 -3582 -3144 -3548
rect -3106 -3582 -3072 -3548
rect -3034 -3582 -3000 -3548
rect -2962 -3582 -2928 -3548
rect -2890 -3582 -2856 -3548
rect -2818 -3582 -2784 -3548
rect -2746 -3582 -2712 -3548
rect -2674 -3582 -2640 -3548
rect -2602 -3582 -2568 -3548
rect -2530 -3582 -2496 -3548
rect -2458 -3582 -2424 -3548
rect -2386 -3582 -2352 -3548
rect -2314 -3582 -2280 -3548
rect -2242 -3582 -2208 -3548
rect -2170 -3582 -2136 -3548
rect -2098 -3582 -2064 -3548
rect -2026 -3582 -1992 -3548
rect -1954 -3582 -1920 -3548
rect -1882 -3582 -1848 -3548
rect -1810 -3582 -1776 -3548
rect -1738 -3582 -1704 -3548
rect -1666 -3582 -1632 -3548
rect -1594 -3582 -1560 -3548
rect -1522 -3582 -1488 -3548
rect -1450 -3582 -1416 -3548
rect -1378 -3582 -1344 -3548
rect -1306 -3582 -1272 -3548
rect -1234 -3582 -1200 -3548
rect -1162 -3582 -1128 -3548
rect -1090 -3582 -1056 -3548
rect -1018 -3582 -984 -3548
rect -946 -3582 -912 -3548
rect -874 -3582 -840 -3548
rect -802 -3582 -768 -3548
rect -730 -3582 -696 -3548
rect -658 -3582 -624 -3548
rect -586 -3582 -552 -3548
rect -514 -3582 -480 -3548
rect -442 -3582 -408 -3548
rect -370 -3582 -336 -3548
rect -298 -3582 -264 -3548
rect -226 -3582 -192 -3548
rect -154 -3582 -120 -3548
rect -82 -3582 -48 -3548
rect -10 -3582 24 -3548
rect 62 -3582 96 -3548
rect 134 -3582 168 -3548
rect 206 -3582 240 -3548
rect 278 -3582 312 -3548
rect 350 -3582 384 -3548
rect 422 -3582 456 -3548
rect 494 -3582 528 -3548
rect 566 -3582 600 -3548
rect 638 -3582 672 -3548
rect 710 -3582 744 -3548
rect 782 -3582 816 -3548
rect 854 -3582 888 -3548
rect 926 -3582 960 -3548
rect 998 -3582 1032 -3548
rect 1070 -3582 1104 -3548
rect 1142 -3582 1176 -3548
rect 1214 -3582 1248 -3548
rect 1286 -3582 1320 -3548
rect 1358 -3582 1392 -3548
rect 1430 -3582 1464 -3548
rect 1502 -3582 1536 -3548
rect 1574 -3582 1608 -3548
rect 1646 -3582 1680 -3548
rect 1718 -3582 1752 -3548
rect 1790 -3582 1824 -3548
rect 1862 -3582 1896 -3548
rect 1934 -3582 1968 -3548
rect 2006 -3582 2040 -3548
rect 2078 -3582 2112 -3548
rect 2150 -3582 2184 -3548
rect 2222 -3582 2256 -3548
rect 2610 -2534 2644 -2500
rect 2610 -2606 2644 -2572
rect 2610 -2678 2644 -2644
rect 2610 -2750 2644 -2716
rect 2610 -2822 2644 -2788
rect 2610 -2894 2644 -2860
rect 2610 -2966 2644 -2932
rect 2610 -3038 2644 -3004
rect 2610 -3110 2644 -3076
rect 2610 -3182 2644 -3148
rect 2576 -3481 2682 -3231
rect -4371 -3730 -4337 -3696
rect -4299 -3730 -4265 -3696
rect -4227 -3730 -4193 -3696
rect -4155 -3730 -4121 -3696
rect -4083 -3730 -4049 -3696
rect -4011 -3730 -3977 -3696
rect -3939 -3730 -3905 -3696
rect -3867 -3730 -3833 -3696
rect -3795 -3730 -3761 -3696
rect -3723 -3730 -3689 -3696
rect -3651 -3730 -3617 -3696
rect -3579 -3730 -3545 -3696
rect -3507 -3730 -3473 -3696
rect -3435 -3730 -3401 -3696
rect -3363 -3730 -3329 -3696
rect -3291 -3730 -3257 -3696
rect -3219 -3730 -3185 -3696
rect -3147 -3730 -3113 -3696
rect -3075 -3730 -3041 -3696
rect -3003 -3730 -2969 -3696
rect -2931 -3730 -2897 -3696
rect -2859 -3730 -2825 -3696
rect -2787 -3730 -2753 -3696
rect -2715 -3730 -2681 -3696
rect -2643 -3730 -2609 -3696
rect -2571 -3730 -2537 -3696
rect -2499 -3730 -2465 -3696
rect -2427 -3730 -2393 -3696
rect -2355 -3730 -2321 -3696
rect -2283 -3730 -2249 -3696
rect -2211 -3730 -2177 -3696
rect -2139 -3730 -2105 -3696
rect -2067 -3730 -2033 -3696
rect -1995 -3730 -1961 -3696
rect -1923 -3730 -1889 -3696
rect -1851 -3730 -1817 -3696
rect -1779 -3730 -1745 -3696
rect -1707 -3730 -1673 -3696
rect -1635 -3730 -1601 -3696
rect -1563 -3730 -1529 -3696
rect -1491 -3730 -1457 -3696
rect -1419 -3730 -1385 -3696
rect -1347 -3730 -1313 -3696
rect -1275 -3730 -1241 -3696
rect -1203 -3730 -1169 -3696
rect -1131 -3730 -1097 -3696
rect -1059 -3730 -1025 -3696
rect -987 -3730 -953 -3696
rect -915 -3730 -881 -3696
rect -843 -3730 -809 -3696
rect -771 -3730 -737 -3696
rect -699 -3730 -665 -3696
rect -627 -3730 -593 -3696
rect -555 -3730 -521 -3696
rect -483 -3730 -449 -3696
rect -411 -3730 -377 -3696
rect -339 -3730 -305 -3696
rect -267 -3730 -233 -3696
rect -195 -3730 -161 -3696
rect -123 -3730 -89 -3696
rect -51 -3730 -17 -3696
rect 21 -3730 55 -3696
rect 93 -3730 127 -3696
rect 165 -3730 199 -3696
rect 237 -3730 271 -3696
rect 309 -3730 343 -3696
rect 381 -3730 415 -3696
rect 453 -3730 487 -3696
rect 525 -3730 559 -3696
rect 597 -3730 631 -3696
rect 669 -3730 703 -3696
rect 741 -3730 775 -3696
rect 813 -3730 847 -3696
rect 885 -3730 919 -3696
rect 957 -3730 991 -3696
rect 1029 -3730 1063 -3696
rect 1101 -3730 1135 -3696
rect 1173 -3730 1207 -3696
rect 1245 -3730 1279 -3696
rect 1317 -3730 1351 -3696
rect 1389 -3730 1423 -3696
rect 1461 -3730 1495 -3696
rect 1533 -3730 1567 -3696
rect 1605 -3730 1639 -3696
rect 1677 -3730 1711 -3696
rect 1749 -3730 1783 -3696
rect 1821 -3730 1855 -3696
rect 1893 -3730 1927 -3696
rect 1965 -3730 1999 -3696
rect 2037 -3730 2071 -3696
rect 2109 -3730 2143 -3696
rect 2181 -3730 2215 -3696
rect 2253 -3730 2287 -3696
rect 2325 -3730 2359 -3696
rect 2397 -3730 2431 -3696
rect 2469 -3730 2503 -3696
rect 2541 -3730 2575 -3696
rect 2613 -3730 2647 -3696
<< metal1 >>
rect -4365 6475 2686 6531
rect -4365 6359 -4326 6475
rect 2638 6359 2686 6475
rect -4365 6316 2686 6359
rect -4365 6296 -4234 6316
rect -4365 6262 -4318 6296
rect -4284 6262 -4234 6296
rect -4365 6224 -4234 6262
rect -4365 6190 -4318 6224
rect -4284 6190 -4234 6224
rect -4365 6152 -4234 6190
rect -4365 6118 -4318 6152
rect -4284 6118 -4234 6152
rect -4365 6080 -4234 6118
rect -4365 6046 -4318 6080
rect -4284 6046 -4234 6080
rect -4365 6008 -4234 6046
rect -4365 5974 -4318 6008
rect -4284 5974 -4234 6008
rect -4365 5936 -4234 5974
rect -4365 5902 -4318 5936
rect -4284 5902 -4234 5936
rect -4365 5864 -4234 5902
rect -4365 5830 -4318 5864
rect -4284 5830 -4234 5864
rect -4365 5792 -4234 5830
rect -4365 5758 -4318 5792
rect -4284 5758 -4234 5792
rect -4365 5720 -4234 5758
rect -4365 5686 -4318 5720
rect -4284 5686 -4234 5720
rect -4365 5648 -4234 5686
rect -4365 5614 -4318 5648
rect -4284 5614 -4234 5648
rect -4365 5576 -4234 5614
rect -4365 5542 -4318 5576
rect -4284 5542 -4234 5576
rect -4365 5504 -4234 5542
rect -4365 5470 -4318 5504
rect -4284 5470 -4234 5504
rect -4365 5432 -4234 5470
rect -4365 5398 -4318 5432
rect -4284 5398 -4234 5432
rect -4365 5360 -4234 5398
rect -4365 5326 -4318 5360
rect -4284 5326 -4234 5360
rect -4365 5288 -4234 5326
rect -4365 5254 -4318 5288
rect -4284 5254 -4234 5288
rect -4365 5216 -4234 5254
rect -4365 5182 -4318 5216
rect -4284 5182 -4234 5216
rect -4365 5144 -4234 5182
rect -4365 5110 -4318 5144
rect -4284 5110 -4234 5144
rect -4365 5072 -4234 5110
rect -4365 5038 -4318 5072
rect -4284 5038 -4234 5072
rect -4365 5000 -4234 5038
rect -4365 4966 -4318 5000
rect -4284 4966 -4234 5000
rect -4365 4928 -4234 4966
rect -4365 4894 -4318 4928
rect -4284 4894 -4234 4928
rect -4365 4856 -4234 4894
rect -4365 4822 -4318 4856
rect -4284 4822 -4234 4856
rect -4365 4784 -4234 4822
rect -4365 4750 -4318 4784
rect -4284 4750 -4234 4784
rect -4365 4712 -4234 4750
rect -4365 4678 -4318 4712
rect -4284 4678 -4234 4712
rect -4365 4640 -4234 4678
rect -4365 4606 -4318 4640
rect -4284 4606 -4234 4640
rect -4365 4568 -4234 4606
rect -4365 4534 -4318 4568
rect -4284 4534 -4234 4568
rect -4365 4496 -4234 4534
rect -4365 4462 -4318 4496
rect -4284 4462 -4234 4496
rect -4365 4424 -4234 4462
rect -4365 4390 -4318 4424
rect -4284 4390 -4234 4424
rect -4365 4352 -4234 4390
rect -4365 4318 -4318 4352
rect -4284 4318 -4234 4352
rect -4365 4280 -4234 4318
rect -4365 4246 -4318 4280
rect -4284 4246 -4234 4280
rect -4365 4208 -4234 4246
rect -4365 4174 -4318 4208
rect -4284 4174 -4234 4208
rect -4365 4140 -4234 4174
rect -4171 6114 2470 6178
rect -4171 5787 -4107 6114
rect -4072 6049 -3944 6055
rect -4072 5997 -4066 6049
rect -4014 5997 -4002 6049
rect -3950 5997 -3944 6049
rect -4072 5991 -3944 5997
rect -3756 6049 -3628 6055
rect -3756 5997 -3750 6049
rect -3698 5997 -3686 6049
rect -3634 5997 -3628 6049
rect -3756 5991 -3628 5997
rect -3440 6049 -3312 6055
rect -3440 5997 -3434 6049
rect -3382 5997 -3370 6049
rect -3318 5997 -3312 6049
rect -3440 5991 -3312 5997
rect -3124 6049 -2996 6055
rect -3124 5997 -3118 6049
rect -3066 5997 -3054 6049
rect -3002 5997 -2996 6049
rect -3124 5991 -2996 5997
rect -2808 6049 -2680 6055
rect -2808 5997 -2802 6049
rect -2750 5997 -2738 6049
rect -2686 5997 -2680 6049
rect -2808 5991 -2680 5997
rect -2492 6049 -2364 6055
rect -2492 5997 -2486 6049
rect -2434 5997 -2422 6049
rect -2370 5997 -2364 6049
rect -2492 5991 -2364 5997
rect -2176 6049 -2048 6055
rect -2176 5997 -2170 6049
rect -2118 5997 -2106 6049
rect -2054 5997 -2048 6049
rect -2176 5991 -2048 5997
rect -1860 6049 -1732 6055
rect -1860 5997 -1854 6049
rect -1802 5997 -1790 6049
rect -1738 5997 -1732 6049
rect -1860 5991 -1732 5997
rect -1544 6049 -1416 6055
rect -1544 5997 -1538 6049
rect -1486 5997 -1474 6049
rect -1422 5997 -1416 6049
rect -1544 5991 -1416 5997
rect -1228 6049 -1100 6055
rect -1228 5997 -1222 6049
rect -1170 5997 -1158 6049
rect -1106 5997 -1100 6049
rect -1228 5991 -1100 5997
rect -912 6049 -784 6055
rect -912 5997 -906 6049
rect -854 5997 -842 6049
rect -790 5997 -784 6049
rect -912 5991 -784 5997
rect -596 6049 -468 6055
rect -596 5997 -590 6049
rect -538 5997 -526 6049
rect -474 5997 -468 6049
rect -596 5991 -468 5997
rect -280 6049 -152 6055
rect -280 5997 -274 6049
rect -222 5997 -210 6049
rect -158 5997 -152 6049
rect -280 5991 -152 5997
rect 36 6049 164 6055
rect 36 5997 42 6049
rect 94 5997 106 6049
rect 158 5997 164 6049
rect 36 5991 164 5997
rect 352 6049 480 6055
rect 352 5997 358 6049
rect 410 5997 422 6049
rect 474 5997 480 6049
rect 352 5991 480 5997
rect 668 6049 796 6055
rect 668 5997 674 6049
rect 726 5997 738 6049
rect 790 5997 796 6049
rect 668 5991 796 5997
rect 984 6049 1112 6055
rect 984 5997 990 6049
rect 1042 5997 1054 6049
rect 1106 5997 1112 6049
rect 984 5991 1112 5997
rect 1300 6049 1428 6055
rect 1300 5997 1306 6049
rect 1358 5997 1370 6049
rect 1422 5997 1428 6049
rect 1300 5991 1428 5997
rect 1616 6049 1744 6055
rect 1616 5997 1622 6049
rect 1674 5997 1686 6049
rect 1738 5997 1744 6049
rect 1616 5991 1744 5997
rect 1932 6049 2060 6055
rect 1932 5997 1938 6049
rect 1990 5997 2002 6049
rect 2054 5997 2060 6049
rect 1932 5991 2060 5997
rect 2248 6049 2376 6055
rect 2248 5997 2254 6049
rect 2306 5997 2318 6049
rect 2370 5997 2376 6049
rect 2248 5991 2376 5997
rect -3914 5924 -3786 5930
rect -3914 5872 -3908 5924
rect -3856 5872 -3844 5924
rect -3792 5872 -3786 5924
rect -3914 5866 -3786 5872
rect -3598 5924 -3470 5930
rect -3598 5872 -3592 5924
rect -3540 5872 -3528 5924
rect -3476 5872 -3470 5924
rect -3598 5866 -3470 5872
rect -3282 5924 -3154 5930
rect -3282 5872 -3276 5924
rect -3224 5872 -3212 5924
rect -3160 5872 -3154 5924
rect -3282 5866 -3154 5872
rect -2966 5924 -2838 5930
rect -2966 5872 -2960 5924
rect -2908 5872 -2896 5924
rect -2844 5872 -2838 5924
rect -2966 5866 -2838 5872
rect -2650 5924 -2522 5930
rect -2650 5872 -2644 5924
rect -2592 5872 -2580 5924
rect -2528 5872 -2522 5924
rect -2650 5866 -2522 5872
rect -2334 5924 -2206 5930
rect -2334 5872 -2328 5924
rect -2276 5872 -2264 5924
rect -2212 5872 -2206 5924
rect -2334 5866 -2206 5872
rect -2018 5924 -1890 5930
rect -2018 5872 -2012 5924
rect -1960 5872 -1948 5924
rect -1896 5872 -1890 5924
rect -2018 5866 -1890 5872
rect -1702 5924 -1574 5930
rect -1702 5872 -1696 5924
rect -1644 5872 -1632 5924
rect -1580 5872 -1574 5924
rect -1702 5866 -1574 5872
rect -1386 5924 -1258 5930
rect -1386 5872 -1380 5924
rect -1328 5872 -1316 5924
rect -1264 5872 -1258 5924
rect -1386 5866 -1258 5872
rect -1070 5924 -942 5930
rect -1070 5872 -1064 5924
rect -1012 5872 -1000 5924
rect -948 5872 -942 5924
rect -1070 5866 -942 5872
rect -754 5924 -626 5930
rect -754 5872 -748 5924
rect -696 5872 -684 5924
rect -632 5872 -626 5924
rect -754 5866 -626 5872
rect -438 5924 -310 5930
rect -438 5872 -432 5924
rect -380 5872 -368 5924
rect -316 5872 -310 5924
rect -438 5866 -310 5872
rect -122 5924 6 5930
rect -122 5872 -116 5924
rect -64 5872 -52 5924
rect 0 5872 6 5924
rect -122 5866 6 5872
rect 194 5924 322 5930
rect 194 5872 200 5924
rect 252 5872 264 5924
rect 316 5872 322 5924
rect 194 5866 322 5872
rect 510 5924 638 5930
rect 510 5872 516 5924
rect 568 5872 580 5924
rect 632 5872 638 5924
rect 510 5866 638 5872
rect 826 5924 954 5930
rect 826 5872 832 5924
rect 884 5872 896 5924
rect 948 5872 954 5924
rect 826 5866 954 5872
rect 1142 5924 1270 5930
rect 1142 5872 1148 5924
rect 1200 5872 1212 5924
rect 1264 5872 1270 5924
rect 1142 5866 1270 5872
rect 1458 5924 1586 5930
rect 1458 5872 1464 5924
rect 1516 5872 1528 5924
rect 1580 5872 1586 5924
rect 1458 5866 1586 5872
rect 1774 5924 1902 5930
rect 1774 5872 1780 5924
rect 1832 5872 1844 5924
rect 1896 5872 1902 5924
rect 1774 5866 1902 5872
rect 2090 5924 2218 5930
rect 2090 5872 2096 5924
rect 2148 5872 2160 5924
rect 2212 5872 2218 5924
rect 2090 5866 2218 5872
rect 2406 5787 2470 6114
rect -4171 5672 2470 5787
rect -4171 5360 -4107 5672
rect -4072 5609 -3944 5615
rect -4072 5557 -4066 5609
rect -4014 5557 -4002 5609
rect -3950 5557 -3944 5609
rect -4072 5551 -3944 5557
rect -3756 5609 -3628 5615
rect -3756 5557 -3750 5609
rect -3698 5557 -3686 5609
rect -3634 5557 -3628 5609
rect -3756 5551 -3628 5557
rect -3440 5609 -3312 5615
rect -3440 5557 -3434 5609
rect -3382 5557 -3370 5609
rect -3318 5557 -3312 5609
rect -3440 5551 -3312 5557
rect -3124 5609 -2996 5615
rect -3124 5557 -3118 5609
rect -3066 5557 -3054 5609
rect -3002 5557 -2996 5609
rect -3124 5551 -2996 5557
rect -2808 5609 -2680 5615
rect -2808 5557 -2802 5609
rect -2750 5557 -2738 5609
rect -2686 5557 -2680 5609
rect -2808 5551 -2680 5557
rect -2492 5609 -2364 5615
rect -2492 5557 -2486 5609
rect -2434 5557 -2422 5609
rect -2370 5557 -2364 5609
rect -2492 5551 -2364 5557
rect -2176 5609 -2048 5615
rect -2176 5557 -2170 5609
rect -2118 5557 -2106 5609
rect -2054 5557 -2048 5609
rect -2176 5551 -2048 5557
rect -1860 5609 -1732 5615
rect -1860 5557 -1854 5609
rect -1802 5557 -1790 5609
rect -1738 5557 -1732 5609
rect -1860 5551 -1732 5557
rect -1544 5609 -1416 5615
rect -1544 5557 -1538 5609
rect -1486 5557 -1474 5609
rect -1422 5557 -1416 5609
rect -1544 5551 -1416 5557
rect -1228 5609 -1100 5615
rect -1228 5557 -1222 5609
rect -1170 5557 -1158 5609
rect -1106 5557 -1100 5609
rect -1228 5551 -1100 5557
rect -912 5609 -784 5615
rect -912 5557 -906 5609
rect -854 5557 -842 5609
rect -790 5557 -784 5609
rect -912 5551 -784 5557
rect -596 5609 -468 5615
rect -596 5557 -590 5609
rect -538 5557 -526 5609
rect -474 5557 -468 5609
rect -596 5551 -468 5557
rect -280 5609 -152 5615
rect -280 5557 -274 5609
rect -222 5557 -210 5609
rect -158 5557 -152 5609
rect -280 5551 -152 5557
rect 36 5609 164 5615
rect 36 5557 42 5609
rect 94 5557 106 5609
rect 158 5557 164 5609
rect 36 5551 164 5557
rect 352 5609 480 5615
rect 352 5557 358 5609
rect 410 5557 422 5609
rect 474 5557 480 5609
rect 352 5551 480 5557
rect 668 5609 796 5615
rect 668 5557 674 5609
rect 726 5557 738 5609
rect 790 5557 796 5609
rect 668 5551 796 5557
rect 984 5609 1112 5615
rect 984 5557 990 5609
rect 1042 5557 1054 5609
rect 1106 5557 1112 5609
rect 984 5551 1112 5557
rect 1300 5609 1428 5615
rect 1300 5557 1306 5609
rect 1358 5557 1370 5609
rect 1422 5557 1428 5609
rect 1300 5551 1428 5557
rect 1616 5609 1744 5615
rect 1616 5557 1622 5609
rect 1674 5557 1686 5609
rect 1738 5557 1744 5609
rect 1616 5551 1744 5557
rect 1932 5609 2060 5615
rect 1932 5557 1938 5609
rect 1990 5557 2002 5609
rect 2054 5557 2060 5609
rect 1932 5551 2060 5557
rect 2248 5609 2376 5615
rect 2248 5557 2254 5609
rect 2306 5557 2318 5609
rect 2370 5557 2376 5609
rect 2248 5551 2376 5557
rect -3914 5484 -3786 5490
rect -3914 5432 -3908 5484
rect -3856 5432 -3844 5484
rect -3792 5432 -3786 5484
rect -3914 5426 -3786 5432
rect -3598 5484 -3470 5490
rect -3598 5432 -3592 5484
rect -3540 5432 -3528 5484
rect -3476 5432 -3470 5484
rect -3598 5426 -3470 5432
rect -3282 5484 -3154 5490
rect -3282 5432 -3276 5484
rect -3224 5432 -3212 5484
rect -3160 5432 -3154 5484
rect -3282 5426 -3154 5432
rect -2966 5484 -2838 5490
rect -2966 5432 -2960 5484
rect -2908 5432 -2896 5484
rect -2844 5432 -2838 5484
rect -2966 5426 -2838 5432
rect -2650 5484 -2522 5490
rect -2650 5432 -2644 5484
rect -2592 5432 -2580 5484
rect -2528 5432 -2522 5484
rect -2650 5426 -2522 5432
rect -2334 5484 -2206 5490
rect -2334 5432 -2328 5484
rect -2276 5432 -2264 5484
rect -2212 5432 -2206 5484
rect -2334 5426 -2206 5432
rect -2018 5484 -1890 5490
rect -2018 5432 -2012 5484
rect -1960 5432 -1948 5484
rect -1896 5432 -1890 5484
rect -2018 5426 -1890 5432
rect -1702 5484 -1574 5490
rect -1702 5432 -1696 5484
rect -1644 5432 -1632 5484
rect -1580 5432 -1574 5484
rect -1702 5426 -1574 5432
rect -1386 5484 -1258 5490
rect -1386 5432 -1380 5484
rect -1328 5432 -1316 5484
rect -1264 5432 -1258 5484
rect -1386 5426 -1258 5432
rect -1070 5484 -942 5490
rect -1070 5432 -1064 5484
rect -1012 5432 -1000 5484
rect -948 5432 -942 5484
rect -1070 5426 -942 5432
rect -754 5484 -626 5490
rect -754 5432 -748 5484
rect -696 5432 -684 5484
rect -632 5432 -626 5484
rect -754 5426 -626 5432
rect -438 5484 -310 5490
rect -438 5432 -432 5484
rect -380 5432 -368 5484
rect -316 5432 -310 5484
rect -438 5426 -310 5432
rect -122 5484 6 5490
rect -122 5432 -116 5484
rect -64 5432 -52 5484
rect 0 5432 6 5484
rect -122 5426 6 5432
rect 194 5484 322 5490
rect 194 5432 200 5484
rect 252 5432 264 5484
rect 316 5432 322 5484
rect 194 5426 322 5432
rect 510 5484 638 5490
rect 510 5432 516 5484
rect 568 5432 580 5484
rect 632 5432 638 5484
rect 510 5426 638 5432
rect 826 5484 954 5490
rect 826 5432 832 5484
rect 884 5432 896 5484
rect 948 5432 954 5484
rect 826 5426 954 5432
rect 1142 5484 1270 5490
rect 1142 5432 1148 5484
rect 1200 5432 1212 5484
rect 1264 5432 1270 5484
rect 1142 5426 1270 5432
rect 1458 5484 1586 5490
rect 1458 5432 1464 5484
rect 1516 5432 1528 5484
rect 1580 5432 1586 5484
rect 1458 5426 1586 5432
rect 1774 5484 1902 5490
rect 1774 5432 1780 5484
rect 1832 5432 1844 5484
rect 1896 5432 1902 5484
rect 1774 5426 1902 5432
rect 2090 5484 2218 5490
rect 2090 5432 2096 5484
rect 2148 5432 2160 5484
rect 2212 5432 2218 5484
rect 2090 5426 2218 5432
rect 2406 5360 2470 5672
rect -4171 5245 2470 5360
rect -4171 4917 -4107 5245
rect -4072 5169 -3944 5175
rect -4072 5117 -4066 5169
rect -4014 5117 -4002 5169
rect -3950 5117 -3944 5169
rect -4072 5111 -3944 5117
rect -3756 5169 -3628 5175
rect -3756 5117 -3750 5169
rect -3698 5117 -3686 5169
rect -3634 5117 -3628 5169
rect -3756 5111 -3628 5117
rect -3440 5169 -3312 5175
rect -3440 5117 -3434 5169
rect -3382 5117 -3370 5169
rect -3318 5117 -3312 5169
rect -3440 5111 -3312 5117
rect -3124 5169 -2996 5175
rect -3124 5117 -3118 5169
rect -3066 5117 -3054 5169
rect -3002 5117 -2996 5169
rect -3124 5111 -2996 5117
rect -2808 5169 -2680 5175
rect -2808 5117 -2802 5169
rect -2750 5117 -2738 5169
rect -2686 5117 -2680 5169
rect -2808 5111 -2680 5117
rect -2492 5169 -2364 5175
rect -2492 5117 -2486 5169
rect -2434 5117 -2422 5169
rect -2370 5117 -2364 5169
rect -2492 5111 -2364 5117
rect -2176 5169 -2048 5175
rect -2176 5117 -2170 5169
rect -2118 5117 -2106 5169
rect -2054 5117 -2048 5169
rect -2176 5111 -2048 5117
rect -1860 5169 -1732 5175
rect -1860 5117 -1854 5169
rect -1802 5117 -1790 5169
rect -1738 5117 -1732 5169
rect -1860 5111 -1732 5117
rect -1544 5169 -1416 5175
rect -1544 5117 -1538 5169
rect -1486 5117 -1474 5169
rect -1422 5117 -1416 5169
rect -1544 5111 -1416 5117
rect -1228 5169 -1100 5175
rect -1228 5117 -1222 5169
rect -1170 5117 -1158 5169
rect -1106 5117 -1100 5169
rect -1228 5111 -1100 5117
rect -912 5169 -784 5175
rect -912 5117 -906 5169
rect -854 5117 -842 5169
rect -790 5117 -784 5169
rect -912 5111 -784 5117
rect -596 5169 -468 5175
rect -596 5117 -590 5169
rect -538 5117 -526 5169
rect -474 5117 -468 5169
rect -596 5111 -468 5117
rect -280 5169 -152 5175
rect -280 5117 -274 5169
rect -222 5117 -210 5169
rect -158 5117 -152 5169
rect -280 5111 -152 5117
rect 36 5169 164 5175
rect 36 5117 42 5169
rect 94 5117 106 5169
rect 158 5117 164 5169
rect 36 5111 164 5117
rect 352 5169 480 5175
rect 352 5117 358 5169
rect 410 5117 422 5169
rect 474 5117 480 5169
rect 352 5111 480 5117
rect 668 5169 796 5175
rect 668 5117 674 5169
rect 726 5117 738 5169
rect 790 5117 796 5169
rect 668 5111 796 5117
rect 984 5169 1112 5175
rect 984 5117 990 5169
rect 1042 5117 1054 5169
rect 1106 5117 1112 5169
rect 984 5111 1112 5117
rect 1300 5169 1428 5175
rect 1300 5117 1306 5169
rect 1358 5117 1370 5169
rect 1422 5117 1428 5169
rect 1300 5111 1428 5117
rect 1616 5169 1744 5175
rect 1616 5117 1622 5169
rect 1674 5117 1686 5169
rect 1738 5117 1744 5169
rect 1616 5111 1744 5117
rect 1932 5169 2060 5175
rect 1932 5117 1938 5169
rect 1990 5117 2002 5169
rect 2054 5117 2060 5169
rect 1932 5111 2060 5117
rect 2248 5169 2376 5175
rect 2248 5117 2254 5169
rect 2306 5117 2318 5169
rect 2370 5117 2376 5169
rect 2248 5111 2376 5117
rect -3914 5044 -3786 5050
rect -3914 4992 -3908 5044
rect -3856 4992 -3844 5044
rect -3792 4992 -3786 5044
rect -3914 4986 -3786 4992
rect -3598 5044 -3470 5050
rect -3598 4992 -3592 5044
rect -3540 4992 -3528 5044
rect -3476 4992 -3470 5044
rect -3598 4986 -3470 4992
rect -3282 5044 -3154 5050
rect -3282 4992 -3276 5044
rect -3224 4992 -3212 5044
rect -3160 4992 -3154 5044
rect -3282 4986 -3154 4992
rect -2966 5044 -2838 5050
rect -2966 4992 -2960 5044
rect -2908 4992 -2896 5044
rect -2844 4992 -2838 5044
rect -2966 4986 -2838 4992
rect -2650 5044 -2522 5050
rect -2650 4992 -2644 5044
rect -2592 4992 -2580 5044
rect -2528 4992 -2522 5044
rect -2650 4986 -2522 4992
rect -2334 5044 -2206 5050
rect -2334 4992 -2328 5044
rect -2276 4992 -2264 5044
rect -2212 4992 -2206 5044
rect -2334 4986 -2206 4992
rect -2018 5044 -1890 5050
rect -2018 4992 -2012 5044
rect -1960 4992 -1948 5044
rect -1896 4992 -1890 5044
rect -2018 4986 -1890 4992
rect -1702 5044 -1574 5050
rect -1702 4992 -1696 5044
rect -1644 4992 -1632 5044
rect -1580 4992 -1574 5044
rect -1702 4986 -1574 4992
rect -1386 5044 -1258 5050
rect -1386 4992 -1380 5044
rect -1328 4992 -1316 5044
rect -1264 4992 -1258 5044
rect -1386 4986 -1258 4992
rect -1070 5044 -942 5050
rect -1070 4992 -1064 5044
rect -1012 4992 -1000 5044
rect -948 4992 -942 5044
rect -1070 4986 -942 4992
rect -754 5044 -626 5050
rect -754 4992 -748 5044
rect -696 4992 -684 5044
rect -632 4992 -626 5044
rect -754 4986 -626 4992
rect -438 5044 -310 5050
rect -438 4992 -432 5044
rect -380 4992 -368 5044
rect -316 4992 -310 5044
rect -438 4986 -310 4992
rect -122 5044 6 5050
rect -122 4992 -116 5044
rect -64 4992 -52 5044
rect 0 4992 6 5044
rect -122 4986 6 4992
rect 194 5044 322 5050
rect 194 4992 200 5044
rect 252 4992 264 5044
rect 316 4992 322 5044
rect 194 4986 322 4992
rect 510 5044 638 5050
rect 510 4992 516 5044
rect 568 4992 580 5044
rect 632 4992 638 5044
rect 510 4986 638 4992
rect 826 5044 954 5050
rect 826 4992 832 5044
rect 884 4992 896 5044
rect 948 4992 954 5044
rect 826 4986 954 4992
rect 1142 5044 1270 5050
rect 1142 4992 1148 5044
rect 1200 4992 1212 5044
rect 1264 4992 1270 5044
rect 1142 4986 1270 4992
rect 1458 5044 1586 5050
rect 1458 4992 1464 5044
rect 1516 4992 1528 5044
rect 1580 4992 1586 5044
rect 1458 4986 1586 4992
rect 1774 5044 1902 5050
rect 1774 4992 1780 5044
rect 1832 4992 1844 5044
rect 1896 4992 1902 5044
rect 1774 4986 1902 4992
rect 2090 5044 2218 5050
rect 2090 4992 2096 5044
rect 2148 4992 2160 5044
rect 2212 4992 2218 5044
rect 2090 4986 2218 4992
rect 2406 4917 2470 5245
rect -4171 4802 2470 4917
rect -4171 4484 -4107 4802
rect -4072 4734 -3944 4740
rect -4072 4682 -4066 4734
rect -4014 4682 -4002 4734
rect -3950 4682 -3944 4734
rect -4072 4676 -3944 4682
rect -3756 4734 -3628 4740
rect -3756 4682 -3750 4734
rect -3698 4682 -3686 4734
rect -3634 4682 -3628 4734
rect -3756 4676 -3628 4682
rect -3440 4734 -3312 4740
rect -3440 4682 -3434 4734
rect -3382 4682 -3370 4734
rect -3318 4682 -3312 4734
rect -3440 4676 -3312 4682
rect -3124 4734 -2996 4740
rect -3124 4682 -3118 4734
rect -3066 4682 -3054 4734
rect -3002 4682 -2996 4734
rect -3124 4676 -2996 4682
rect -2808 4734 -2680 4740
rect -2808 4682 -2802 4734
rect -2750 4682 -2738 4734
rect -2686 4682 -2680 4734
rect -2808 4676 -2680 4682
rect -2492 4734 -2364 4740
rect -2492 4682 -2486 4734
rect -2434 4682 -2422 4734
rect -2370 4682 -2364 4734
rect -2492 4676 -2364 4682
rect -2176 4734 -2048 4740
rect -2176 4682 -2170 4734
rect -2118 4682 -2106 4734
rect -2054 4682 -2048 4734
rect -2176 4676 -2048 4682
rect -1860 4734 -1732 4740
rect -1860 4682 -1854 4734
rect -1802 4682 -1790 4734
rect -1738 4682 -1732 4734
rect -1860 4676 -1732 4682
rect -1544 4734 -1416 4740
rect -1544 4682 -1538 4734
rect -1486 4682 -1474 4734
rect -1422 4682 -1416 4734
rect -1544 4676 -1416 4682
rect -1228 4734 -1100 4740
rect -1228 4682 -1222 4734
rect -1170 4682 -1158 4734
rect -1106 4682 -1100 4734
rect -1228 4676 -1100 4682
rect -912 4734 -784 4740
rect -912 4682 -906 4734
rect -854 4682 -842 4734
rect -790 4682 -784 4734
rect -912 4676 -784 4682
rect -596 4734 -468 4740
rect -596 4682 -590 4734
rect -538 4682 -526 4734
rect -474 4682 -468 4734
rect -596 4676 -468 4682
rect -280 4734 -152 4740
rect -280 4682 -274 4734
rect -222 4682 -210 4734
rect -158 4682 -152 4734
rect -280 4676 -152 4682
rect 36 4734 164 4740
rect 36 4682 42 4734
rect 94 4682 106 4734
rect 158 4682 164 4734
rect 36 4676 164 4682
rect 352 4734 480 4740
rect 352 4682 358 4734
rect 410 4682 422 4734
rect 474 4682 480 4734
rect 352 4676 480 4682
rect 668 4734 796 4740
rect 668 4682 674 4734
rect 726 4682 738 4734
rect 790 4682 796 4734
rect 668 4676 796 4682
rect 984 4734 1112 4740
rect 984 4682 990 4734
rect 1042 4682 1054 4734
rect 1106 4682 1112 4734
rect 984 4676 1112 4682
rect 1300 4734 1428 4740
rect 1300 4682 1306 4734
rect 1358 4682 1370 4734
rect 1422 4682 1428 4734
rect 1300 4676 1428 4682
rect 1616 4734 1744 4740
rect 1616 4682 1622 4734
rect 1674 4682 1686 4734
rect 1738 4682 1744 4734
rect 1616 4676 1744 4682
rect 1932 4734 2060 4740
rect 1932 4682 1938 4734
rect 1990 4682 2002 4734
rect 2054 4682 2060 4734
rect 1932 4676 2060 4682
rect 2248 4734 2376 4740
rect 2248 4682 2254 4734
rect 2306 4682 2318 4734
rect 2370 4682 2376 4734
rect 2248 4676 2376 4682
rect -3914 4609 -3786 4615
rect -3914 4557 -3908 4609
rect -3856 4557 -3844 4609
rect -3792 4557 -3786 4609
rect -3914 4551 -3786 4557
rect -3598 4609 -3470 4615
rect -3598 4557 -3592 4609
rect -3540 4557 -3528 4609
rect -3476 4557 -3470 4609
rect -3598 4551 -3470 4557
rect -3282 4609 -3154 4615
rect -3282 4557 -3276 4609
rect -3224 4557 -3212 4609
rect -3160 4557 -3154 4609
rect -3282 4551 -3154 4557
rect -2966 4609 -2838 4615
rect -2966 4557 -2960 4609
rect -2908 4557 -2896 4609
rect -2844 4557 -2838 4609
rect -2966 4551 -2838 4557
rect -2650 4609 -2522 4615
rect -2650 4557 -2644 4609
rect -2592 4557 -2580 4609
rect -2528 4557 -2522 4609
rect -2650 4551 -2522 4557
rect -2334 4609 -2206 4615
rect -2334 4557 -2328 4609
rect -2276 4557 -2264 4609
rect -2212 4557 -2206 4609
rect -2334 4551 -2206 4557
rect -2018 4609 -1890 4615
rect -2018 4557 -2012 4609
rect -1960 4557 -1948 4609
rect -1896 4557 -1890 4609
rect -2018 4551 -1890 4557
rect -1702 4609 -1574 4615
rect -1702 4557 -1696 4609
rect -1644 4557 -1632 4609
rect -1580 4557 -1574 4609
rect -1702 4551 -1574 4557
rect -1386 4609 -1258 4615
rect -1386 4557 -1380 4609
rect -1328 4557 -1316 4609
rect -1264 4557 -1258 4609
rect -1386 4551 -1258 4557
rect -1070 4609 -942 4615
rect -1070 4557 -1064 4609
rect -1012 4557 -1000 4609
rect -948 4557 -942 4609
rect -1070 4551 -942 4557
rect -754 4609 -626 4615
rect -754 4557 -748 4609
rect -696 4557 -684 4609
rect -632 4557 -626 4609
rect -754 4551 -626 4557
rect -438 4609 -310 4615
rect -438 4557 -432 4609
rect -380 4557 -368 4609
rect -316 4557 -310 4609
rect -438 4551 -310 4557
rect -122 4609 6 4615
rect -122 4557 -116 4609
rect -64 4557 -52 4609
rect 0 4557 6 4609
rect -122 4551 6 4557
rect 194 4609 322 4615
rect 194 4557 200 4609
rect 252 4557 264 4609
rect 316 4557 322 4609
rect 194 4551 322 4557
rect 510 4609 638 4615
rect 510 4557 516 4609
rect 568 4557 580 4609
rect 632 4557 638 4609
rect 510 4551 638 4557
rect 826 4609 954 4615
rect 826 4557 832 4609
rect 884 4557 896 4609
rect 948 4557 954 4609
rect 826 4551 954 4557
rect 1142 4609 1270 4615
rect 1142 4557 1148 4609
rect 1200 4557 1212 4609
rect 1264 4557 1270 4609
rect 1142 4551 1270 4557
rect 1458 4609 1586 4615
rect 1458 4557 1464 4609
rect 1516 4557 1528 4609
rect 1580 4557 1586 4609
rect 1458 4551 1586 4557
rect 1774 4609 1902 4615
rect 1774 4557 1780 4609
rect 1832 4557 1844 4609
rect 1896 4557 1902 4609
rect 1774 4551 1902 4557
rect 2090 4609 2218 4615
rect 2090 4557 2096 4609
rect 2148 4557 2160 4609
rect 2212 4557 2218 4609
rect 2090 4551 2218 4557
rect 2406 4484 2470 4802
rect -4171 4369 2470 4484
rect -4171 4071 -4107 4369
rect -4072 4309 -3944 4315
rect -4072 4257 -4066 4309
rect -4014 4257 -4002 4309
rect -3950 4257 -3944 4309
rect -4072 4251 -3944 4257
rect -3756 4309 -3628 4315
rect -3756 4257 -3750 4309
rect -3698 4257 -3686 4309
rect -3634 4257 -3628 4309
rect -3756 4251 -3628 4257
rect -3440 4309 -3312 4315
rect -3440 4257 -3434 4309
rect -3382 4257 -3370 4309
rect -3318 4257 -3312 4309
rect -3440 4251 -3312 4257
rect -3124 4309 -2996 4315
rect -3124 4257 -3118 4309
rect -3066 4257 -3054 4309
rect -3002 4257 -2996 4309
rect -3124 4251 -2996 4257
rect -2808 4309 -2680 4315
rect -2808 4257 -2802 4309
rect -2750 4257 -2738 4309
rect -2686 4257 -2680 4309
rect -2808 4251 -2680 4257
rect -2492 4309 -2364 4315
rect -2492 4257 -2486 4309
rect -2434 4257 -2422 4309
rect -2370 4257 -2364 4309
rect -2492 4251 -2364 4257
rect -2176 4309 -2048 4315
rect -2176 4257 -2170 4309
rect -2118 4257 -2106 4309
rect -2054 4257 -2048 4309
rect -2176 4251 -2048 4257
rect -1860 4309 -1732 4315
rect -1860 4257 -1854 4309
rect -1802 4257 -1790 4309
rect -1738 4257 -1732 4309
rect -1860 4251 -1732 4257
rect -1544 4309 -1416 4315
rect -1544 4257 -1538 4309
rect -1486 4257 -1474 4309
rect -1422 4257 -1416 4309
rect -1544 4251 -1416 4257
rect -1228 4309 -1100 4315
rect -1228 4257 -1222 4309
rect -1170 4257 -1158 4309
rect -1106 4257 -1100 4309
rect -1228 4251 -1100 4257
rect -912 4309 -784 4315
rect -912 4257 -906 4309
rect -854 4257 -842 4309
rect -790 4257 -784 4309
rect -912 4251 -784 4257
rect -596 4309 -468 4315
rect -596 4257 -590 4309
rect -538 4257 -526 4309
rect -474 4257 -468 4309
rect -596 4251 -468 4257
rect -280 4309 -152 4315
rect -280 4257 -274 4309
rect -222 4257 -210 4309
rect -158 4257 -152 4309
rect -280 4251 -152 4257
rect 36 4309 164 4315
rect 36 4257 42 4309
rect 94 4257 106 4309
rect 158 4257 164 4309
rect 36 4251 164 4257
rect 352 4309 480 4315
rect 352 4257 358 4309
rect 410 4257 422 4309
rect 474 4257 480 4309
rect 352 4251 480 4257
rect 668 4309 796 4315
rect 668 4257 674 4309
rect 726 4257 738 4309
rect 790 4257 796 4309
rect 668 4251 796 4257
rect 984 4309 1112 4315
rect 984 4257 990 4309
rect 1042 4257 1054 4309
rect 1106 4257 1112 4309
rect 984 4251 1112 4257
rect 1300 4309 1428 4315
rect 1300 4257 1306 4309
rect 1358 4257 1370 4309
rect 1422 4257 1428 4309
rect 1300 4251 1428 4257
rect 1616 4309 1744 4315
rect 1616 4257 1622 4309
rect 1674 4257 1686 4309
rect 1738 4257 1744 4309
rect 1616 4251 1744 4257
rect 1932 4309 2060 4315
rect 1932 4257 1938 4309
rect 1990 4257 2002 4309
rect 2054 4257 2060 4309
rect 1932 4251 2060 4257
rect 2248 4309 2376 4315
rect 2248 4257 2254 4309
rect 2306 4257 2318 4309
rect 2370 4257 2376 4309
rect 2248 4251 2376 4257
rect -3914 4184 -3786 4190
rect -3914 4132 -3908 4184
rect -3856 4132 -3844 4184
rect -3792 4132 -3786 4184
rect -3914 4126 -3786 4132
rect -3598 4184 -3470 4190
rect -3598 4132 -3592 4184
rect -3540 4132 -3528 4184
rect -3476 4132 -3470 4184
rect -3598 4126 -3470 4132
rect -3282 4184 -3154 4190
rect -3282 4132 -3276 4184
rect -3224 4132 -3212 4184
rect -3160 4132 -3154 4184
rect -3282 4126 -3154 4132
rect -2966 4184 -2838 4190
rect -2966 4132 -2960 4184
rect -2908 4132 -2896 4184
rect -2844 4132 -2838 4184
rect -2966 4126 -2838 4132
rect -2650 4184 -2522 4190
rect -2650 4132 -2644 4184
rect -2592 4132 -2580 4184
rect -2528 4132 -2522 4184
rect -2650 4126 -2522 4132
rect -2334 4184 -2206 4190
rect -2334 4132 -2328 4184
rect -2276 4132 -2264 4184
rect -2212 4132 -2206 4184
rect -2334 4126 -2206 4132
rect -2018 4184 -1890 4190
rect -2018 4132 -2012 4184
rect -1960 4132 -1948 4184
rect -1896 4132 -1890 4184
rect -2018 4126 -1890 4132
rect -1702 4184 -1574 4190
rect -1702 4132 -1696 4184
rect -1644 4132 -1632 4184
rect -1580 4132 -1574 4184
rect -1702 4126 -1574 4132
rect -1386 4184 -1258 4190
rect -1386 4132 -1380 4184
rect -1328 4132 -1316 4184
rect -1264 4132 -1258 4184
rect -1386 4126 -1258 4132
rect -1070 4184 -942 4190
rect -1070 4132 -1064 4184
rect -1012 4132 -1000 4184
rect -948 4132 -942 4184
rect -1070 4126 -942 4132
rect -754 4184 -626 4190
rect -754 4132 -748 4184
rect -696 4132 -684 4184
rect -632 4132 -626 4184
rect -754 4126 -626 4132
rect -438 4184 -310 4190
rect -438 4132 -432 4184
rect -380 4132 -368 4184
rect -316 4132 -310 4184
rect -438 4126 -310 4132
rect -122 4184 6 4190
rect -122 4132 -116 4184
rect -64 4132 -52 4184
rect 0 4132 6 4184
rect -122 4126 6 4132
rect 194 4184 322 4190
rect 194 4132 200 4184
rect 252 4132 264 4184
rect 316 4132 322 4184
rect 194 4126 322 4132
rect 510 4184 638 4190
rect 510 4132 516 4184
rect 568 4132 580 4184
rect 632 4132 638 4184
rect 510 4126 638 4132
rect 826 4184 954 4190
rect 826 4132 832 4184
rect 884 4132 896 4184
rect 948 4132 954 4184
rect 826 4126 954 4132
rect 1142 4184 1270 4190
rect 1142 4132 1148 4184
rect 1200 4132 1212 4184
rect 1264 4132 1270 4184
rect 1142 4126 1270 4132
rect 1458 4184 1586 4190
rect 1458 4132 1464 4184
rect 1516 4132 1528 4184
rect 1580 4132 1586 4184
rect 1458 4126 1586 4132
rect 1774 4184 1902 4190
rect 1774 4132 1780 4184
rect 1832 4132 1844 4184
rect 1896 4132 1902 4184
rect 1774 4126 1902 4132
rect 2090 4184 2218 4190
rect 2090 4132 2096 4184
rect 2148 4132 2160 4184
rect 2212 4132 2218 4184
rect 2090 4126 2218 4132
rect -4291 4066 -4107 4071
rect 2406 4066 2470 4369
rect -4291 4002 2470 4066
rect 2534 6104 2683 6131
rect -4291 1583 -4227 4002
rect -4170 3937 2485 3941
rect -4170 3926 -4110 3937
rect -4058 3926 -4046 3937
rect -3994 3926 -3982 3937
rect -3930 3926 -3918 3937
rect -3866 3926 -3854 3937
rect -4170 3892 -4148 3926
rect -4114 3892 -4110 3926
rect -3866 3892 -3860 3926
rect -4170 3885 -4110 3892
rect -4058 3885 -4046 3892
rect -3994 3885 -3982 3892
rect -3930 3885 -3918 3892
rect -3866 3885 -3854 3892
rect -3802 3885 -3790 3937
rect -3738 3885 -3726 3937
rect -3674 3885 -3662 3937
rect -3610 3885 -3598 3937
rect -3546 3926 -3534 3937
rect -3482 3926 -3470 3937
rect -3418 3926 -3406 3937
rect -3354 3926 -3342 3937
rect -3290 3926 -3278 3937
rect -3538 3892 -3534 3926
rect -3290 3892 -3284 3926
rect -3546 3885 -3534 3892
rect -3482 3885 -3470 3892
rect -3418 3885 -3406 3892
rect -3354 3885 -3342 3892
rect -3290 3885 -3278 3892
rect -3226 3885 -3214 3937
rect -3162 3885 -3150 3937
rect -3098 3885 -3086 3937
rect -3034 3885 -3022 3937
rect -2970 3926 -2958 3937
rect -2906 3926 -2894 3937
rect -2842 3926 -2830 3937
rect -2778 3926 -2766 3937
rect -2714 3926 -2702 3937
rect -2962 3892 -2958 3926
rect -2714 3892 -2708 3926
rect -2970 3885 -2958 3892
rect -2906 3885 -2894 3892
rect -2842 3885 -2830 3892
rect -2778 3885 -2766 3892
rect -2714 3885 -2702 3892
rect -2650 3885 -2638 3937
rect -2586 3885 -2574 3937
rect -2522 3885 -2510 3937
rect -2458 3885 -2446 3937
rect -2394 3926 -2382 3937
rect -2330 3926 -2318 3937
rect -2266 3926 -2254 3937
rect -2202 3926 -2190 3937
rect -2138 3926 -2126 3937
rect -2386 3892 -2382 3926
rect -2138 3892 -2132 3926
rect -2394 3885 -2382 3892
rect -2330 3885 -2318 3892
rect -2266 3885 -2254 3892
rect -2202 3885 -2190 3892
rect -2138 3885 -2126 3892
rect -2074 3885 -2062 3937
rect -2010 3885 -1998 3937
rect -1946 3885 -1934 3937
rect -1882 3885 -1870 3937
rect -1818 3926 -1806 3937
rect -1754 3926 -1742 3937
rect -1690 3926 -1678 3937
rect -1626 3926 -1614 3937
rect -1562 3926 -1550 3937
rect -1810 3892 -1806 3926
rect -1562 3892 -1556 3926
rect -1818 3885 -1806 3892
rect -1754 3885 -1742 3892
rect -1690 3885 -1678 3892
rect -1626 3885 -1614 3892
rect -1562 3885 -1550 3892
rect -1498 3885 -1486 3937
rect -1434 3885 -1422 3937
rect -1370 3885 -1358 3937
rect -1306 3885 -1294 3937
rect -1242 3926 -1230 3937
rect -1178 3926 -1166 3937
rect -1114 3926 -1102 3937
rect -1050 3926 -1038 3937
rect -986 3926 -974 3937
rect -1234 3892 -1230 3926
rect -986 3892 -980 3926
rect -1242 3885 -1230 3892
rect -1178 3885 -1166 3892
rect -1114 3885 -1102 3892
rect -1050 3885 -1038 3892
rect -986 3885 -974 3892
rect -922 3885 -910 3937
rect -858 3885 -846 3937
rect -794 3885 -782 3937
rect -730 3885 -718 3937
rect -666 3926 -654 3937
rect -602 3926 -590 3937
rect -538 3926 -526 3937
rect -474 3926 -462 3937
rect -410 3926 -398 3937
rect -658 3892 -654 3926
rect -410 3892 -404 3926
rect -666 3885 -654 3892
rect -602 3885 -590 3892
rect -538 3885 -526 3892
rect -474 3885 -462 3892
rect -410 3885 -398 3892
rect -346 3885 -334 3937
rect -282 3885 -270 3937
rect -218 3885 -206 3937
rect -154 3885 -142 3937
rect -90 3926 -78 3937
rect -26 3926 -14 3937
rect 38 3926 50 3937
rect 102 3926 114 3937
rect 166 3926 178 3937
rect -82 3892 -78 3926
rect 166 3892 172 3926
rect -90 3885 -78 3892
rect -26 3885 -14 3892
rect 38 3885 50 3892
rect 102 3885 114 3892
rect 166 3885 178 3892
rect 230 3885 242 3937
rect 294 3885 306 3937
rect 358 3885 370 3937
rect 422 3885 434 3937
rect 486 3926 498 3937
rect 550 3926 562 3937
rect 614 3926 626 3937
rect 678 3926 690 3937
rect 742 3926 754 3937
rect 494 3892 498 3926
rect 742 3892 748 3926
rect 486 3885 498 3892
rect 550 3885 562 3892
rect 614 3885 626 3892
rect 678 3885 690 3892
rect 742 3885 754 3892
rect 806 3885 818 3937
rect 870 3885 882 3937
rect 934 3885 946 3937
rect 998 3885 1010 3937
rect 1062 3926 1074 3937
rect 1126 3926 1138 3937
rect 1190 3926 1202 3937
rect 1254 3926 1266 3937
rect 1318 3926 1330 3937
rect 1070 3892 1074 3926
rect 1318 3892 1324 3926
rect 1062 3885 1074 3892
rect 1126 3885 1138 3892
rect 1190 3885 1202 3892
rect 1254 3885 1266 3892
rect 1318 3885 1330 3892
rect 1382 3885 1394 3937
rect 1446 3885 1458 3937
rect 1510 3885 1522 3937
rect 1574 3885 1586 3937
rect 1638 3926 1650 3937
rect 1702 3926 1714 3937
rect 1766 3926 1778 3937
rect 1830 3926 1842 3937
rect 1894 3926 1906 3937
rect 1646 3892 1650 3926
rect 1894 3892 1900 3926
rect 1638 3885 1650 3892
rect 1702 3885 1714 3892
rect 1766 3885 1778 3892
rect 1830 3885 1842 3892
rect 1894 3885 1906 3892
rect 1958 3885 1970 3937
rect 2022 3885 2034 3937
rect 2086 3885 2098 3937
rect 2150 3885 2162 3937
rect 2214 3926 2226 3937
rect 2278 3926 2290 3937
rect 2342 3926 2485 3937
rect 2222 3892 2226 3926
rect 2366 3892 2404 3926
rect 2438 3892 2485 3926
rect 2214 3885 2226 3892
rect 2278 3885 2290 3892
rect 2342 3885 2485 3892
rect -4170 3881 2485 3885
rect -4174 3757 2476 3821
rect -4174 3440 -4110 3757
rect -4072 3689 -3944 3695
rect -4072 3637 -4066 3689
rect -4014 3637 -4002 3689
rect -3950 3637 -3944 3689
rect -4072 3631 -3944 3637
rect -3756 3689 -3628 3695
rect -3756 3637 -3750 3689
rect -3698 3637 -3686 3689
rect -3634 3637 -3628 3689
rect -3756 3631 -3628 3637
rect -3440 3689 -3312 3695
rect -3440 3637 -3434 3689
rect -3382 3637 -3370 3689
rect -3318 3637 -3312 3689
rect -3440 3631 -3312 3637
rect -3124 3689 -2996 3695
rect -3124 3637 -3118 3689
rect -3066 3637 -3054 3689
rect -3002 3637 -2996 3689
rect -3124 3631 -2996 3637
rect -2808 3689 -2680 3695
rect -2808 3637 -2802 3689
rect -2750 3637 -2738 3689
rect -2686 3637 -2680 3689
rect -2808 3631 -2680 3637
rect -2492 3689 -2364 3695
rect -2492 3637 -2486 3689
rect -2434 3637 -2422 3689
rect -2370 3637 -2364 3689
rect -2492 3631 -2364 3637
rect -2176 3689 -2048 3695
rect -2176 3637 -2170 3689
rect -2118 3637 -2106 3689
rect -2054 3637 -2048 3689
rect -2176 3631 -2048 3637
rect -1860 3689 -1732 3695
rect -1860 3637 -1854 3689
rect -1802 3637 -1790 3689
rect -1738 3637 -1732 3689
rect -1860 3631 -1732 3637
rect -1544 3689 -1416 3695
rect -1544 3637 -1538 3689
rect -1486 3637 -1474 3689
rect -1422 3637 -1416 3689
rect -1544 3631 -1416 3637
rect -1228 3689 -1100 3695
rect -1228 3637 -1222 3689
rect -1170 3637 -1158 3689
rect -1106 3637 -1100 3689
rect -1228 3631 -1100 3637
rect -912 3689 -784 3695
rect -912 3637 -906 3689
rect -854 3637 -842 3689
rect -790 3637 -784 3689
rect -912 3631 -784 3637
rect -596 3689 -468 3695
rect -596 3637 -590 3689
rect -538 3637 -526 3689
rect -474 3637 -468 3689
rect -596 3631 -468 3637
rect -280 3689 -152 3695
rect -280 3637 -274 3689
rect -222 3637 -210 3689
rect -158 3637 -152 3689
rect -280 3631 -152 3637
rect 36 3689 164 3695
rect 36 3637 42 3689
rect 94 3637 106 3689
rect 158 3637 164 3689
rect 36 3631 164 3637
rect 352 3689 480 3695
rect 352 3637 358 3689
rect 410 3637 422 3689
rect 474 3637 480 3689
rect 352 3631 480 3637
rect 668 3689 796 3695
rect 668 3637 674 3689
rect 726 3637 738 3689
rect 790 3637 796 3689
rect 668 3631 796 3637
rect 984 3689 1112 3695
rect 984 3637 990 3689
rect 1042 3637 1054 3689
rect 1106 3637 1112 3689
rect 984 3631 1112 3637
rect 1300 3689 1428 3695
rect 1300 3637 1306 3689
rect 1358 3637 1370 3689
rect 1422 3637 1428 3689
rect 1300 3631 1428 3637
rect 1616 3689 1744 3695
rect 1616 3637 1622 3689
rect 1674 3637 1686 3689
rect 1738 3637 1744 3689
rect 1616 3631 1744 3637
rect 1932 3689 2060 3695
rect 1932 3637 1938 3689
rect 1990 3637 2002 3689
rect 2054 3637 2060 3689
rect 1932 3631 2060 3637
rect 2248 3689 2376 3695
rect 2248 3637 2254 3689
rect 2306 3637 2318 3689
rect 2370 3637 2376 3689
rect 2248 3631 2376 3637
rect -3914 3564 -3786 3570
rect -3914 3512 -3908 3564
rect -3856 3512 -3844 3564
rect -3792 3512 -3786 3564
rect -3914 3506 -3786 3512
rect -3598 3564 -3470 3570
rect -3598 3512 -3592 3564
rect -3540 3512 -3528 3564
rect -3476 3512 -3470 3564
rect -3598 3506 -3470 3512
rect -3282 3564 -3154 3570
rect -3282 3512 -3276 3564
rect -3224 3512 -3212 3564
rect -3160 3512 -3154 3564
rect -3282 3506 -3154 3512
rect -2966 3564 -2838 3570
rect -2966 3512 -2960 3564
rect -2908 3512 -2896 3564
rect -2844 3512 -2838 3564
rect -2966 3506 -2838 3512
rect -2650 3564 -2522 3570
rect -2650 3512 -2644 3564
rect -2592 3512 -2580 3564
rect -2528 3512 -2522 3564
rect -2650 3506 -2522 3512
rect -2334 3564 -2206 3570
rect -2334 3512 -2328 3564
rect -2276 3512 -2264 3564
rect -2212 3512 -2206 3564
rect -2334 3506 -2206 3512
rect -2018 3564 -1890 3570
rect -2018 3512 -2012 3564
rect -1960 3512 -1948 3564
rect -1896 3512 -1890 3564
rect -2018 3506 -1890 3512
rect -1702 3564 -1574 3570
rect -1702 3512 -1696 3564
rect -1644 3512 -1632 3564
rect -1580 3512 -1574 3564
rect -1702 3506 -1574 3512
rect -1386 3564 -1258 3570
rect -1386 3512 -1380 3564
rect -1328 3512 -1316 3564
rect -1264 3512 -1258 3564
rect -1386 3506 -1258 3512
rect -1070 3564 -942 3570
rect -1070 3512 -1064 3564
rect -1012 3512 -1000 3564
rect -948 3512 -942 3564
rect -1070 3506 -942 3512
rect -754 3564 -626 3570
rect -754 3512 -748 3564
rect -696 3512 -684 3564
rect -632 3512 -626 3564
rect -754 3506 -626 3512
rect -438 3564 -310 3570
rect -438 3512 -432 3564
rect -380 3512 -368 3564
rect -316 3512 -310 3564
rect -438 3506 -310 3512
rect -122 3564 6 3570
rect -122 3512 -116 3564
rect -64 3512 -52 3564
rect 0 3512 6 3564
rect -122 3506 6 3512
rect 194 3564 322 3570
rect 194 3512 200 3564
rect 252 3512 264 3564
rect 316 3512 322 3564
rect 194 3506 322 3512
rect 510 3564 638 3570
rect 510 3512 516 3564
rect 568 3512 580 3564
rect 632 3512 638 3564
rect 510 3506 638 3512
rect 826 3564 954 3570
rect 826 3512 832 3564
rect 884 3512 896 3564
rect 948 3512 954 3564
rect 826 3506 954 3512
rect 1142 3564 1270 3570
rect 1142 3512 1148 3564
rect 1200 3512 1212 3564
rect 1264 3512 1270 3564
rect 1142 3506 1270 3512
rect 1458 3564 1586 3570
rect 1458 3512 1464 3564
rect 1516 3512 1528 3564
rect 1580 3512 1586 3564
rect 1458 3506 1586 3512
rect 1774 3564 1902 3570
rect 1774 3512 1780 3564
rect 1832 3512 1844 3564
rect 1896 3512 1902 3564
rect 1774 3506 1902 3512
rect 2090 3564 2218 3570
rect 2090 3512 2096 3564
rect 2148 3512 2160 3564
rect 2212 3512 2218 3564
rect 2090 3506 2218 3512
rect 2412 3440 2476 3757
rect -4174 3325 2476 3440
rect -4174 3002 -4110 3325
rect -4072 3254 -3944 3260
rect -4072 3202 -4066 3254
rect -4014 3202 -4002 3254
rect -3950 3202 -3944 3254
rect -4072 3196 -3944 3202
rect -3756 3254 -3628 3260
rect -3756 3202 -3750 3254
rect -3698 3202 -3686 3254
rect -3634 3202 -3628 3254
rect -3756 3196 -3628 3202
rect -3440 3254 -3312 3260
rect -3440 3202 -3434 3254
rect -3382 3202 -3370 3254
rect -3318 3202 -3312 3254
rect -3440 3196 -3312 3202
rect -3124 3254 -2996 3260
rect -3124 3202 -3118 3254
rect -3066 3202 -3054 3254
rect -3002 3202 -2996 3254
rect -3124 3196 -2996 3202
rect -2808 3254 -2680 3260
rect -2808 3202 -2802 3254
rect -2750 3202 -2738 3254
rect -2686 3202 -2680 3254
rect -2808 3196 -2680 3202
rect -2492 3254 -2364 3260
rect -2492 3202 -2486 3254
rect -2434 3202 -2422 3254
rect -2370 3202 -2364 3254
rect -2492 3196 -2364 3202
rect -2176 3254 -2048 3260
rect -2176 3202 -2170 3254
rect -2118 3202 -2106 3254
rect -2054 3202 -2048 3254
rect -2176 3196 -2048 3202
rect -1860 3254 -1732 3260
rect -1860 3202 -1854 3254
rect -1802 3202 -1790 3254
rect -1738 3202 -1732 3254
rect -1860 3196 -1732 3202
rect -1544 3254 -1416 3260
rect -1544 3202 -1538 3254
rect -1486 3202 -1474 3254
rect -1422 3202 -1416 3254
rect -1544 3196 -1416 3202
rect -1228 3254 -1100 3260
rect -1228 3202 -1222 3254
rect -1170 3202 -1158 3254
rect -1106 3202 -1100 3254
rect -1228 3196 -1100 3202
rect -912 3254 -784 3260
rect -912 3202 -906 3254
rect -854 3202 -842 3254
rect -790 3202 -784 3254
rect -912 3196 -784 3202
rect -596 3254 -468 3260
rect -596 3202 -590 3254
rect -538 3202 -526 3254
rect -474 3202 -468 3254
rect -596 3196 -468 3202
rect -280 3254 -152 3260
rect -280 3202 -274 3254
rect -222 3202 -210 3254
rect -158 3202 -152 3254
rect -280 3196 -152 3202
rect 36 3254 164 3260
rect 36 3202 42 3254
rect 94 3202 106 3254
rect 158 3202 164 3254
rect 36 3196 164 3202
rect 352 3254 480 3260
rect 352 3202 358 3254
rect 410 3202 422 3254
rect 474 3202 480 3254
rect 352 3196 480 3202
rect 668 3254 796 3260
rect 668 3202 674 3254
rect 726 3202 738 3254
rect 790 3202 796 3254
rect 668 3196 796 3202
rect 984 3254 1112 3260
rect 984 3202 990 3254
rect 1042 3202 1054 3254
rect 1106 3202 1112 3254
rect 984 3196 1112 3202
rect 1300 3254 1428 3260
rect 1300 3202 1306 3254
rect 1358 3202 1370 3254
rect 1422 3202 1428 3254
rect 1300 3196 1428 3202
rect 1616 3254 1744 3260
rect 1616 3202 1622 3254
rect 1674 3202 1686 3254
rect 1738 3202 1744 3254
rect 1616 3196 1744 3202
rect 1932 3254 2060 3260
rect 1932 3202 1938 3254
rect 1990 3202 2002 3254
rect 2054 3202 2060 3254
rect 1932 3196 2060 3202
rect 2248 3254 2376 3260
rect 2248 3202 2254 3254
rect 2306 3202 2318 3254
rect 2370 3202 2376 3254
rect 2248 3196 2376 3202
rect -3914 3129 -3786 3135
rect -3914 3077 -3908 3129
rect -3856 3077 -3844 3129
rect -3792 3077 -3786 3129
rect -3914 3071 -3786 3077
rect -3598 3129 -3470 3135
rect -3598 3077 -3592 3129
rect -3540 3077 -3528 3129
rect -3476 3077 -3470 3129
rect -3598 3071 -3470 3077
rect -3282 3129 -3154 3135
rect -3282 3077 -3276 3129
rect -3224 3077 -3212 3129
rect -3160 3077 -3154 3129
rect -3282 3071 -3154 3077
rect -2966 3129 -2838 3135
rect -2966 3077 -2960 3129
rect -2908 3077 -2896 3129
rect -2844 3077 -2838 3129
rect -2966 3071 -2838 3077
rect -2650 3129 -2522 3135
rect -2650 3077 -2644 3129
rect -2592 3077 -2580 3129
rect -2528 3077 -2522 3129
rect -2650 3071 -2522 3077
rect -2334 3129 -2206 3135
rect -2334 3077 -2328 3129
rect -2276 3077 -2264 3129
rect -2212 3077 -2206 3129
rect -2334 3071 -2206 3077
rect -2018 3129 -1890 3135
rect -2018 3077 -2012 3129
rect -1960 3077 -1948 3129
rect -1896 3077 -1890 3129
rect -2018 3071 -1890 3077
rect -1702 3129 -1574 3135
rect -1702 3077 -1696 3129
rect -1644 3077 -1632 3129
rect -1580 3077 -1574 3129
rect -1702 3071 -1574 3077
rect -1386 3129 -1258 3135
rect -1386 3077 -1380 3129
rect -1328 3077 -1316 3129
rect -1264 3077 -1258 3129
rect -1386 3071 -1258 3077
rect -1070 3129 -942 3135
rect -1070 3077 -1064 3129
rect -1012 3077 -1000 3129
rect -948 3077 -942 3129
rect -1070 3071 -942 3077
rect -754 3129 -626 3135
rect -754 3077 -748 3129
rect -696 3077 -684 3129
rect -632 3077 -626 3129
rect -754 3071 -626 3077
rect -438 3129 -310 3135
rect -438 3077 -432 3129
rect -380 3077 -368 3129
rect -316 3077 -310 3129
rect -438 3071 -310 3077
rect -122 3129 6 3135
rect -122 3077 -116 3129
rect -64 3077 -52 3129
rect 0 3077 6 3129
rect -122 3071 6 3077
rect 194 3129 322 3135
rect 194 3077 200 3129
rect 252 3077 264 3129
rect 316 3077 322 3129
rect 194 3071 322 3077
rect 510 3129 638 3135
rect 510 3077 516 3129
rect 568 3077 580 3129
rect 632 3077 638 3129
rect 510 3071 638 3077
rect 826 3129 954 3135
rect 826 3077 832 3129
rect 884 3077 896 3129
rect 948 3077 954 3129
rect 826 3071 954 3077
rect 1142 3129 1270 3135
rect 1142 3077 1148 3129
rect 1200 3077 1212 3129
rect 1264 3077 1270 3129
rect 1142 3071 1270 3077
rect 1458 3129 1586 3135
rect 1458 3077 1464 3129
rect 1516 3077 1528 3129
rect 1580 3077 1586 3129
rect 1458 3071 1586 3077
rect 1774 3129 1902 3135
rect 1774 3077 1780 3129
rect 1832 3077 1844 3129
rect 1896 3077 1902 3129
rect 1774 3071 1902 3077
rect 2090 3129 2218 3135
rect 2090 3077 2096 3129
rect 2148 3077 2160 3129
rect 2212 3077 2218 3129
rect 2090 3071 2218 3077
rect 2412 3002 2476 3325
rect -4174 2887 2476 3002
rect -4174 2570 -4110 2887
rect -4072 2819 -3944 2825
rect -4072 2767 -4066 2819
rect -4014 2767 -4002 2819
rect -3950 2767 -3944 2819
rect -4072 2761 -3944 2767
rect -3756 2819 -3628 2825
rect -3756 2767 -3750 2819
rect -3698 2767 -3686 2819
rect -3634 2767 -3628 2819
rect -3756 2761 -3628 2767
rect -3440 2819 -3312 2825
rect -3440 2767 -3434 2819
rect -3382 2767 -3370 2819
rect -3318 2767 -3312 2819
rect -3440 2761 -3312 2767
rect -3124 2819 -2996 2825
rect -3124 2767 -3118 2819
rect -3066 2767 -3054 2819
rect -3002 2767 -2996 2819
rect -3124 2761 -2996 2767
rect -2808 2819 -2680 2825
rect -2808 2767 -2802 2819
rect -2750 2767 -2738 2819
rect -2686 2767 -2680 2819
rect -2808 2761 -2680 2767
rect -2492 2819 -2364 2825
rect -2492 2767 -2486 2819
rect -2434 2767 -2422 2819
rect -2370 2767 -2364 2819
rect -2492 2761 -2364 2767
rect -2176 2819 -2048 2825
rect -2176 2767 -2170 2819
rect -2118 2767 -2106 2819
rect -2054 2767 -2048 2819
rect -2176 2761 -2048 2767
rect -1860 2819 -1732 2825
rect -1860 2767 -1854 2819
rect -1802 2767 -1790 2819
rect -1738 2767 -1732 2819
rect -1860 2761 -1732 2767
rect -1544 2819 -1416 2825
rect -1544 2767 -1538 2819
rect -1486 2767 -1474 2819
rect -1422 2767 -1416 2819
rect -1544 2761 -1416 2767
rect -1228 2819 -1100 2825
rect -1228 2767 -1222 2819
rect -1170 2767 -1158 2819
rect -1106 2767 -1100 2819
rect -1228 2761 -1100 2767
rect -912 2819 -784 2825
rect -912 2767 -906 2819
rect -854 2767 -842 2819
rect -790 2767 -784 2819
rect -912 2761 -784 2767
rect -596 2819 -468 2825
rect -596 2767 -590 2819
rect -538 2767 -526 2819
rect -474 2767 -468 2819
rect -596 2761 -468 2767
rect -280 2819 -152 2825
rect -280 2767 -274 2819
rect -222 2767 -210 2819
rect -158 2767 -152 2819
rect -280 2761 -152 2767
rect 36 2819 164 2825
rect 36 2767 42 2819
rect 94 2767 106 2819
rect 158 2767 164 2819
rect 36 2761 164 2767
rect 352 2819 480 2825
rect 352 2767 358 2819
rect 410 2767 422 2819
rect 474 2767 480 2819
rect 352 2761 480 2767
rect 668 2819 796 2825
rect 668 2767 674 2819
rect 726 2767 738 2819
rect 790 2767 796 2819
rect 668 2761 796 2767
rect 984 2819 1112 2825
rect 984 2767 990 2819
rect 1042 2767 1054 2819
rect 1106 2767 1112 2819
rect 984 2761 1112 2767
rect 1300 2819 1428 2825
rect 1300 2767 1306 2819
rect 1358 2767 1370 2819
rect 1422 2767 1428 2819
rect 1300 2761 1428 2767
rect 1616 2819 1744 2825
rect 1616 2767 1622 2819
rect 1674 2767 1686 2819
rect 1738 2767 1744 2819
rect 1616 2761 1744 2767
rect 1932 2819 2060 2825
rect 1932 2767 1938 2819
rect 1990 2767 2002 2819
rect 2054 2767 2060 2819
rect 1932 2761 2060 2767
rect 2248 2819 2376 2825
rect 2248 2767 2254 2819
rect 2306 2767 2318 2819
rect 2370 2767 2376 2819
rect 2248 2761 2376 2767
rect -3914 2694 -3786 2700
rect -3914 2642 -3908 2694
rect -3856 2642 -3844 2694
rect -3792 2642 -3786 2694
rect -3914 2636 -3786 2642
rect -3598 2694 -3470 2700
rect -3598 2642 -3592 2694
rect -3540 2642 -3528 2694
rect -3476 2642 -3470 2694
rect -3598 2636 -3470 2642
rect -3282 2694 -3154 2700
rect -3282 2642 -3276 2694
rect -3224 2642 -3212 2694
rect -3160 2642 -3154 2694
rect -3282 2636 -3154 2642
rect -2966 2694 -2838 2700
rect -2966 2642 -2960 2694
rect -2908 2642 -2896 2694
rect -2844 2642 -2838 2694
rect -2966 2636 -2838 2642
rect -2650 2694 -2522 2700
rect -2650 2642 -2644 2694
rect -2592 2642 -2580 2694
rect -2528 2642 -2522 2694
rect -2650 2636 -2522 2642
rect -2334 2694 -2206 2700
rect -2334 2642 -2328 2694
rect -2276 2642 -2264 2694
rect -2212 2642 -2206 2694
rect -2334 2636 -2206 2642
rect -2018 2694 -1890 2700
rect -2018 2642 -2012 2694
rect -1960 2642 -1948 2694
rect -1896 2642 -1890 2694
rect -2018 2636 -1890 2642
rect -1702 2694 -1574 2700
rect -1702 2642 -1696 2694
rect -1644 2642 -1632 2694
rect -1580 2642 -1574 2694
rect -1702 2636 -1574 2642
rect -1386 2694 -1258 2700
rect -1386 2642 -1380 2694
rect -1328 2642 -1316 2694
rect -1264 2642 -1258 2694
rect -1386 2636 -1258 2642
rect -1070 2694 -942 2700
rect -1070 2642 -1064 2694
rect -1012 2642 -1000 2694
rect -948 2642 -942 2694
rect -1070 2636 -942 2642
rect -754 2694 -626 2700
rect -754 2642 -748 2694
rect -696 2642 -684 2694
rect -632 2642 -626 2694
rect -754 2636 -626 2642
rect -438 2694 -310 2700
rect -438 2642 -432 2694
rect -380 2642 -368 2694
rect -316 2642 -310 2694
rect -438 2636 -310 2642
rect -122 2694 6 2700
rect -122 2642 -116 2694
rect -64 2642 -52 2694
rect 0 2642 6 2694
rect -122 2636 6 2642
rect 194 2694 322 2700
rect 194 2642 200 2694
rect 252 2642 264 2694
rect 316 2642 322 2694
rect 194 2636 322 2642
rect 510 2694 638 2700
rect 510 2642 516 2694
rect 568 2642 580 2694
rect 632 2642 638 2694
rect 510 2636 638 2642
rect 826 2694 954 2700
rect 826 2642 832 2694
rect 884 2642 896 2694
rect 948 2642 954 2694
rect 826 2636 954 2642
rect 1142 2694 1270 2700
rect 1142 2642 1148 2694
rect 1200 2642 1212 2694
rect 1264 2642 1270 2694
rect 1142 2636 1270 2642
rect 1458 2694 1586 2700
rect 1458 2642 1464 2694
rect 1516 2642 1528 2694
rect 1580 2642 1586 2694
rect 1458 2636 1586 2642
rect 1774 2694 1902 2700
rect 1774 2642 1780 2694
rect 1832 2642 1844 2694
rect 1896 2642 1902 2694
rect 1774 2636 1902 2642
rect 2090 2694 2218 2700
rect 2090 2642 2096 2694
rect 2148 2642 2160 2694
rect 2212 2642 2218 2694
rect 2090 2636 2218 2642
rect 2412 2570 2476 2887
rect -4174 2455 2476 2570
rect -4174 2135 -4110 2455
rect -4072 2384 -3944 2390
rect -4072 2332 -4066 2384
rect -4014 2332 -4002 2384
rect -3950 2332 -3944 2384
rect -4072 2326 -3944 2332
rect -3756 2384 -3628 2390
rect -3756 2332 -3750 2384
rect -3698 2332 -3686 2384
rect -3634 2332 -3628 2384
rect -3756 2326 -3628 2332
rect -3440 2384 -3312 2390
rect -3440 2332 -3434 2384
rect -3382 2332 -3370 2384
rect -3318 2332 -3312 2384
rect -3440 2326 -3312 2332
rect -3124 2384 -2996 2390
rect -3124 2332 -3118 2384
rect -3066 2332 -3054 2384
rect -3002 2332 -2996 2384
rect -3124 2326 -2996 2332
rect -2808 2384 -2680 2390
rect -2808 2332 -2802 2384
rect -2750 2332 -2738 2384
rect -2686 2332 -2680 2384
rect -2808 2326 -2680 2332
rect -2492 2384 -2364 2390
rect -2492 2332 -2486 2384
rect -2434 2332 -2422 2384
rect -2370 2332 -2364 2384
rect -2492 2326 -2364 2332
rect -2176 2384 -2048 2390
rect -2176 2332 -2170 2384
rect -2118 2332 -2106 2384
rect -2054 2332 -2048 2384
rect -2176 2326 -2048 2332
rect -1860 2384 -1732 2390
rect -1860 2332 -1854 2384
rect -1802 2332 -1790 2384
rect -1738 2332 -1732 2384
rect -1860 2326 -1732 2332
rect -1544 2384 -1416 2390
rect -1544 2332 -1538 2384
rect -1486 2332 -1474 2384
rect -1422 2332 -1416 2384
rect -1544 2326 -1416 2332
rect -1228 2384 -1100 2390
rect -1228 2332 -1222 2384
rect -1170 2332 -1158 2384
rect -1106 2332 -1100 2384
rect -1228 2326 -1100 2332
rect -912 2384 -784 2390
rect -912 2332 -906 2384
rect -854 2332 -842 2384
rect -790 2332 -784 2384
rect -912 2326 -784 2332
rect -596 2384 -468 2390
rect -596 2332 -590 2384
rect -538 2332 -526 2384
rect -474 2332 -468 2384
rect -596 2326 -468 2332
rect -280 2384 -152 2390
rect -280 2332 -274 2384
rect -222 2332 -210 2384
rect -158 2332 -152 2384
rect -280 2326 -152 2332
rect 36 2384 164 2390
rect 36 2332 42 2384
rect 94 2332 106 2384
rect 158 2332 164 2384
rect 36 2326 164 2332
rect 352 2384 480 2390
rect 352 2332 358 2384
rect 410 2332 422 2384
rect 474 2332 480 2384
rect 352 2326 480 2332
rect 668 2384 796 2390
rect 668 2332 674 2384
rect 726 2332 738 2384
rect 790 2332 796 2384
rect 668 2326 796 2332
rect 984 2384 1112 2390
rect 984 2332 990 2384
rect 1042 2332 1054 2384
rect 1106 2332 1112 2384
rect 984 2326 1112 2332
rect 1300 2384 1428 2390
rect 1300 2332 1306 2384
rect 1358 2332 1370 2384
rect 1422 2332 1428 2384
rect 1300 2326 1428 2332
rect 1616 2384 1744 2390
rect 1616 2332 1622 2384
rect 1674 2332 1686 2384
rect 1738 2332 1744 2384
rect 1616 2326 1744 2332
rect 1932 2384 2060 2390
rect 1932 2332 1938 2384
rect 1990 2332 2002 2384
rect 2054 2332 2060 2384
rect 1932 2326 2060 2332
rect 2248 2384 2376 2390
rect 2248 2332 2254 2384
rect 2306 2332 2318 2384
rect 2370 2332 2376 2384
rect 2248 2326 2376 2332
rect -3914 2259 -3786 2265
rect -3914 2207 -3908 2259
rect -3856 2207 -3844 2259
rect -3792 2207 -3786 2259
rect -3914 2201 -3786 2207
rect -3598 2259 -3470 2265
rect -3598 2207 -3592 2259
rect -3540 2207 -3528 2259
rect -3476 2207 -3470 2259
rect -3598 2201 -3470 2207
rect -3282 2259 -3154 2265
rect -3282 2207 -3276 2259
rect -3224 2207 -3212 2259
rect -3160 2207 -3154 2259
rect -3282 2201 -3154 2207
rect -2966 2259 -2838 2265
rect -2966 2207 -2960 2259
rect -2908 2207 -2896 2259
rect -2844 2207 -2838 2259
rect -2966 2201 -2838 2207
rect -2650 2259 -2522 2265
rect -2650 2207 -2644 2259
rect -2592 2207 -2580 2259
rect -2528 2207 -2522 2259
rect -2650 2201 -2522 2207
rect -2334 2259 -2206 2265
rect -2334 2207 -2328 2259
rect -2276 2207 -2264 2259
rect -2212 2207 -2206 2259
rect -2334 2201 -2206 2207
rect -2018 2259 -1890 2265
rect -2018 2207 -2012 2259
rect -1960 2207 -1948 2259
rect -1896 2207 -1890 2259
rect -2018 2201 -1890 2207
rect -1702 2259 -1574 2265
rect -1702 2207 -1696 2259
rect -1644 2207 -1632 2259
rect -1580 2207 -1574 2259
rect -1702 2201 -1574 2207
rect -1386 2259 -1258 2265
rect -1386 2207 -1380 2259
rect -1328 2207 -1316 2259
rect -1264 2207 -1258 2259
rect -1386 2201 -1258 2207
rect -1070 2259 -942 2265
rect -1070 2207 -1064 2259
rect -1012 2207 -1000 2259
rect -948 2207 -942 2259
rect -1070 2201 -942 2207
rect -754 2259 -626 2265
rect -754 2207 -748 2259
rect -696 2207 -684 2259
rect -632 2207 -626 2259
rect -754 2201 -626 2207
rect -438 2259 -310 2265
rect -438 2207 -432 2259
rect -380 2207 -368 2259
rect -316 2207 -310 2259
rect -438 2201 -310 2207
rect -122 2259 6 2265
rect -122 2207 -116 2259
rect -64 2207 -52 2259
rect 0 2207 6 2259
rect -122 2201 6 2207
rect 194 2259 322 2265
rect 194 2207 200 2259
rect 252 2207 264 2259
rect 316 2207 322 2259
rect 194 2201 322 2207
rect 510 2259 638 2265
rect 510 2207 516 2259
rect 568 2207 580 2259
rect 632 2207 638 2259
rect 510 2201 638 2207
rect 826 2259 954 2265
rect 826 2207 832 2259
rect 884 2207 896 2259
rect 948 2207 954 2259
rect 826 2201 954 2207
rect 1142 2259 1270 2265
rect 1142 2207 1148 2259
rect 1200 2207 1212 2259
rect 1264 2207 1270 2259
rect 1142 2201 1270 2207
rect 1458 2259 1586 2265
rect 1458 2207 1464 2259
rect 1516 2207 1528 2259
rect 1580 2207 1586 2259
rect 1458 2201 1586 2207
rect 1774 2259 1902 2265
rect 1774 2207 1780 2259
rect 1832 2207 1844 2259
rect 1896 2207 1902 2259
rect 1774 2201 1902 2207
rect 2090 2259 2218 2265
rect 2090 2207 2096 2259
rect 2148 2207 2160 2259
rect 2212 2207 2218 2259
rect 2090 2201 2218 2207
rect 2412 2135 2476 2455
rect -4174 2040 2476 2135
rect -4174 1713 -4110 2040
rect -4072 1949 -3944 1955
rect -4072 1897 -4066 1949
rect -4014 1897 -4002 1949
rect -3950 1897 -3944 1949
rect -4072 1891 -3944 1897
rect -3756 1949 -3628 1955
rect -3756 1897 -3750 1949
rect -3698 1897 -3686 1949
rect -3634 1897 -3628 1949
rect -3756 1891 -3628 1897
rect -3440 1949 -3312 1955
rect -3440 1897 -3434 1949
rect -3382 1897 -3370 1949
rect -3318 1897 -3312 1949
rect -3440 1891 -3312 1897
rect -3124 1949 -2996 1955
rect -3124 1897 -3118 1949
rect -3066 1897 -3054 1949
rect -3002 1897 -2996 1949
rect -3124 1891 -2996 1897
rect -2808 1949 -2680 1955
rect -2808 1897 -2802 1949
rect -2750 1897 -2738 1949
rect -2686 1897 -2680 1949
rect -2808 1891 -2680 1897
rect -2492 1949 -2364 1955
rect -2492 1897 -2486 1949
rect -2434 1897 -2422 1949
rect -2370 1897 -2364 1949
rect -2492 1891 -2364 1897
rect -2176 1949 -2048 1955
rect -2176 1897 -2170 1949
rect -2118 1897 -2106 1949
rect -2054 1897 -2048 1949
rect -2176 1891 -2048 1897
rect -1860 1949 -1732 1955
rect -1860 1897 -1854 1949
rect -1802 1897 -1790 1949
rect -1738 1897 -1732 1949
rect -1860 1891 -1732 1897
rect -1544 1949 -1416 1955
rect -1544 1897 -1538 1949
rect -1486 1897 -1474 1949
rect -1422 1897 -1416 1949
rect -1544 1891 -1416 1897
rect -1228 1949 -1100 1955
rect -1228 1897 -1222 1949
rect -1170 1897 -1158 1949
rect -1106 1897 -1100 1949
rect -1228 1891 -1100 1897
rect -912 1949 -784 1955
rect -912 1897 -906 1949
rect -854 1897 -842 1949
rect -790 1897 -784 1949
rect -912 1891 -784 1897
rect -596 1949 -468 1955
rect -596 1897 -590 1949
rect -538 1897 -526 1949
rect -474 1897 -468 1949
rect -596 1891 -468 1897
rect -280 1949 -152 1955
rect -280 1897 -274 1949
rect -222 1897 -210 1949
rect -158 1897 -152 1949
rect -280 1891 -152 1897
rect 36 1949 164 1955
rect 36 1897 42 1949
rect 94 1897 106 1949
rect 158 1897 164 1949
rect 36 1891 164 1897
rect 352 1949 480 1955
rect 352 1897 358 1949
rect 410 1897 422 1949
rect 474 1897 480 1949
rect 352 1891 480 1897
rect 668 1949 796 1955
rect 668 1897 674 1949
rect 726 1897 738 1949
rect 790 1897 796 1949
rect 668 1891 796 1897
rect 984 1949 1112 1955
rect 984 1897 990 1949
rect 1042 1897 1054 1949
rect 1106 1897 1112 1949
rect 984 1891 1112 1897
rect 1300 1949 1428 1955
rect 1300 1897 1306 1949
rect 1358 1897 1370 1949
rect 1422 1897 1428 1949
rect 1300 1891 1428 1897
rect 1616 1949 1744 1955
rect 1616 1897 1622 1949
rect 1674 1897 1686 1949
rect 1738 1897 1744 1949
rect 1616 1891 1744 1897
rect 1932 1949 2060 1955
rect 1932 1897 1938 1949
rect 1990 1897 2002 1949
rect 2054 1897 2060 1949
rect 1932 1891 2060 1897
rect 2248 1949 2376 1955
rect 2248 1897 2254 1949
rect 2306 1897 2318 1949
rect 2370 1897 2376 1949
rect 2248 1891 2376 1897
rect -3914 1824 -3786 1830
rect -3914 1772 -3908 1824
rect -3856 1772 -3844 1824
rect -3792 1772 -3786 1824
rect -3914 1766 -3786 1772
rect -3598 1824 -3470 1830
rect -3598 1772 -3592 1824
rect -3540 1772 -3528 1824
rect -3476 1772 -3470 1824
rect -3598 1766 -3470 1772
rect -3282 1824 -3154 1830
rect -3282 1772 -3276 1824
rect -3224 1772 -3212 1824
rect -3160 1772 -3154 1824
rect -3282 1766 -3154 1772
rect -2966 1824 -2838 1830
rect -2966 1772 -2960 1824
rect -2908 1772 -2896 1824
rect -2844 1772 -2838 1824
rect -2966 1766 -2838 1772
rect -2650 1824 -2522 1830
rect -2650 1772 -2644 1824
rect -2592 1772 -2580 1824
rect -2528 1772 -2522 1824
rect -2650 1766 -2522 1772
rect -2334 1824 -2206 1830
rect -2334 1772 -2328 1824
rect -2276 1772 -2264 1824
rect -2212 1772 -2206 1824
rect -2334 1766 -2206 1772
rect -2018 1824 -1890 1830
rect -2018 1772 -2012 1824
rect -1960 1772 -1948 1824
rect -1896 1772 -1890 1824
rect -2018 1766 -1890 1772
rect -1702 1824 -1574 1830
rect -1702 1772 -1696 1824
rect -1644 1772 -1632 1824
rect -1580 1772 -1574 1824
rect -1702 1766 -1574 1772
rect -1386 1824 -1258 1830
rect -1386 1772 -1380 1824
rect -1328 1772 -1316 1824
rect -1264 1772 -1258 1824
rect -1386 1766 -1258 1772
rect -1070 1824 -942 1830
rect -1070 1772 -1064 1824
rect -1012 1772 -1000 1824
rect -948 1772 -942 1824
rect -1070 1766 -942 1772
rect -754 1824 -626 1830
rect -754 1772 -748 1824
rect -696 1772 -684 1824
rect -632 1772 -626 1824
rect -754 1766 -626 1772
rect -438 1824 -310 1830
rect -438 1772 -432 1824
rect -380 1772 -368 1824
rect -316 1772 -310 1824
rect -438 1766 -310 1772
rect -122 1824 6 1830
rect -122 1772 -116 1824
rect -64 1772 -52 1824
rect 0 1772 6 1824
rect -122 1766 6 1772
rect 194 1824 322 1830
rect 194 1772 200 1824
rect 252 1772 264 1824
rect 316 1772 322 1824
rect 194 1766 322 1772
rect 510 1824 638 1830
rect 510 1772 516 1824
rect 568 1772 580 1824
rect 632 1772 638 1824
rect 510 1766 638 1772
rect 826 1824 954 1830
rect 826 1772 832 1824
rect 884 1772 896 1824
rect 948 1772 954 1824
rect 826 1766 954 1772
rect 1142 1824 1270 1830
rect 1142 1772 1148 1824
rect 1200 1772 1212 1824
rect 1264 1772 1270 1824
rect 1142 1766 1270 1772
rect 1458 1824 1586 1830
rect 1458 1772 1464 1824
rect 1516 1772 1528 1824
rect 1580 1772 1586 1824
rect 1458 1766 1586 1772
rect 1774 1824 1902 1830
rect 1774 1772 1780 1824
rect 1832 1772 1844 1824
rect 1896 1772 1902 1824
rect 1774 1766 1902 1772
rect 2090 1824 2218 1830
rect 2090 1772 2096 1824
rect 2148 1772 2160 1824
rect 2212 1772 2218 1824
rect 2090 1766 2218 1772
rect 2412 1713 2476 2040
rect -4174 1649 2476 1713
rect -4291 1519 -3634 1583
rect 2412 1569 2476 1649
rect -4362 1179 -4140 1401
rect -4362 1176 -4342 1179
rect -4164 1176 -4140 1179
rect -4077 1400 -3813 1445
rect -4077 1220 -4036 1400
rect -3856 1220 -3813 1400
rect -4077 1177 -3813 1220
rect -4362 932 -4343 1176
rect -4163 932 -4140 1176
rect -4362 929 -4342 932
rect -4164 929 -4140 932
rect -4362 911 -4140 929
rect -4361 779 -3762 789
rect -4361 599 -4098 779
rect -3854 599 -3762 779
rect -4361 589 -3762 599
rect -3846 452 -3762 589
rect -3698 491 -3634 1519
rect 1911 1506 2476 1569
rect 2534 1508 2550 6104
rect 2666 1508 2683 6104
rect 1911 1505 2412 1506
rect -3444 1401 1553 1449
rect -3444 1381 -3173 1401
rect -3444 555 -3397 1381
rect -3291 1366 -3173 1381
rect 1295 1400 1553 1401
rect 1295 1366 1404 1400
rect -3291 1260 -3193 1366
rect 1305 1260 1404 1366
rect -3291 1221 -3173 1260
rect 1295 1221 1404 1260
rect -3291 1181 1404 1221
rect -3291 555 -3246 1181
rect -2947 1177 -1099 1181
rect 447 1177 749 1181
rect -3444 498 -3246 555
rect -3113 596 -3064 840
rect -2947 640 -2854 1177
rect -2746 874 -2386 911
rect -2746 596 -2697 874
rect -3113 560 -2697 596
rect -3113 506 -3064 560
rect -2746 506 -2697 560
rect -2529 507 -2480 840
rect -2423 595 -2386 874
rect -2356 638 -2263 1177
rect -2424 559 -2217 595
rect -2159 507 -2110 840
rect -3705 489 -3522 491
rect -4361 325 -4126 444
rect -3705 437 -3672 489
rect -3620 437 -3608 489
rect -3556 437 -3522 489
rect -3705 436 -3522 437
rect -3113 424 -2697 506
rect -2595 489 -2110 507
rect -2595 437 -2507 489
rect -2455 437 -2443 489
rect -2391 437 -2379 489
rect -2327 437 -2315 489
rect -2263 437 -2251 489
rect -2199 437 -2187 489
rect -2135 437 -2110 489
rect -3113 423 -2701 424
rect -4361 244 -3762 325
rect -3846 213 -3762 244
rect -3228 227 -3210 279
rect -3158 227 -3146 279
rect -3094 227 -3075 279
rect -3846 161 -3828 213
rect -3776 161 -3762 213
rect -3846 149 -3762 161
rect -3846 97 -3828 149
rect -3776 97 -3762 149
rect -4392 15 -3980 34
rect -4392 1 -4105 15
rect -4392 -307 -4344 1
rect -4164 -307 -4105 1
rect -4392 -523 -4105 -307
rect -3999 -198 -3980 15
rect -3846 -143 -3762 97
rect -3537 15 -3380 56
rect -3537 -198 -3509 15
rect -3999 -335 -3509 -198
rect -3999 -523 -3980 -335
rect -3909 -413 -3702 -408
rect -3909 -465 -3861 -413
rect -3809 -465 -3797 -413
rect -3745 -465 -3702 -413
rect -3909 -469 -3702 -465
rect -3537 -451 -3509 -335
rect -3403 -451 -3380 15
rect -3221 -70 -3156 -60
rect -3221 -122 -3214 -70
rect -3162 -122 -3156 -70
rect -3221 -134 -3156 -122
rect -3221 -186 -3214 -134
rect -3162 -186 -3156 -134
rect -3221 -198 -3156 -186
rect -3221 -250 -3214 -198
rect -3162 -250 -3156 -198
rect -3221 -256 -3156 -250
rect -3123 -329 -3084 227
rect -3028 -253 -2937 423
rect -2595 421 -2110 437
rect -1946 595 -1897 840
rect -1779 636 -1686 1177
rect -1578 878 -1220 915
rect -1578 595 -1529 878
rect -1946 559 -1529 595
rect -1946 504 -1897 559
rect -1578 504 -1529 559
rect -1946 423 -1529 504
rect -1356 504 -1307 840
rect -1257 595 -1220 878
rect -1192 638 -1099 1177
rect -1263 559 -1056 595
rect -996 504 -947 840
rect -1356 487 -947 504
rect -1356 435 -1338 487
rect -1286 435 -1274 487
rect -1222 435 -1210 487
rect -1158 435 -1146 487
rect -1094 435 -1082 487
rect -1030 435 -1018 487
rect -966 435 -947 487
rect -2795 323 -2777 375
rect -2725 323 -2713 375
rect -2661 323 -2642 375
rect -2788 -70 -2723 -60
rect -2788 -122 -2776 -70
rect -2724 -122 -2723 -70
rect -2788 -134 -2723 -122
rect -2788 -186 -2776 -134
rect -2724 -186 -2723 -134
rect -2788 -198 -2723 -186
rect -2788 -250 -2776 -198
rect -2724 -250 -2723 -198
rect -2788 -256 -2723 -250
rect -2693 -322 -2653 323
rect -2595 -256 -2505 421
rect -1927 227 -1909 279
rect -1857 227 -1845 279
rect -1793 227 -1774 279
rect -2284 80 -2192 86
rect -2284 28 -2264 80
rect -2212 28 -2192 80
rect -2284 20 -2192 28
rect -4392 -546 -3980 -523
rect -4392 -547 -4120 -546
rect -4434 -667 -4296 -607
rect -3892 -621 -3825 -469
rect -3537 -486 -3380 -451
rect -2407 -531 -2312 -58
rect -2256 -316 -2214 20
rect -2183 -67 -2118 -60
rect -2183 -119 -2178 -67
rect -2126 -119 -2118 -67
rect -2183 -131 -2118 -119
rect -2183 -183 -2178 -131
rect -2126 -183 -2118 -131
rect -2183 -195 -2118 -183
rect -2183 -247 -2178 -195
rect -2126 -247 -2118 -195
rect -2183 -256 -2118 -247
rect -1916 -68 -1851 -60
rect -1916 -120 -1907 -68
rect -1855 -120 -1851 -68
rect -1916 -132 -1851 -120
rect -1916 -184 -1907 -132
rect -1855 -184 -1851 -132
rect -1916 -196 -1851 -184
rect -1916 -248 -1907 -196
rect -1855 -248 -1851 -196
rect -1916 -256 -1851 -248
rect -1822 -329 -1781 227
rect -1724 -253 -1639 423
rect -1356 422 -947 435
rect -1495 323 -1477 375
rect -1425 323 -1413 375
rect -1361 323 -1342 375
rect -1485 -67 -1420 -60
rect -1485 -119 -1478 -67
rect -1426 -119 -1420 -67
rect -1485 -131 -1420 -119
rect -1485 -183 -1478 -131
rect -1426 -183 -1420 -131
rect -1485 -195 -1420 -183
rect -1485 -247 -1478 -195
rect -1426 -247 -1420 -195
rect -1485 -256 -1420 -247
rect -1389 -320 -1350 323
rect -1290 -256 -1199 422
rect -779 153 -733 840
rect -622 832 -510 848
rect -622 780 -592 832
rect -540 780 -510 832
rect -622 768 -510 780
rect -622 716 -592 768
rect -540 716 -510 768
rect -622 704 -510 716
rect -622 652 -592 704
rect -540 652 -510 704
rect -622 638 -510 652
rect -665 375 -624 585
rect -502 375 -461 581
rect -665 323 -654 375
rect -602 323 -590 375
rect -538 323 -526 375
rect -474 323 -461 375
rect -410 153 -364 840
rect -981 80 -889 86
rect -981 28 -961 80
rect -909 28 -889 80
rect -779 54 -364 153
rect -191 152 -145 840
rect -36 830 76 847
rect -36 778 -7 830
rect 45 778 76 830
rect -36 766 76 778
rect -36 714 -7 766
rect 45 714 76 766
rect -36 702 76 714
rect -36 650 -7 702
rect 45 650 76 702
rect -36 637 76 650
rect -85 279 -44 580
rect 74 279 115 582
rect -86 227 -75 279
rect -23 227 -11 279
rect 41 227 53 279
rect 105 227 116 279
rect 185 152 231 840
rect 388 830 500 846
rect 388 778 415 830
rect 467 778 500 830
rect 388 766 500 778
rect 388 714 415 766
rect 467 714 500 766
rect 388 702 500 714
rect 388 650 415 702
rect 467 650 500 702
rect 388 636 500 650
rect 539 640 667 1177
rect 707 833 819 849
rect 707 781 735 833
rect 787 781 819 833
rect 707 769 819 781
rect 707 717 735 769
rect 787 717 819 769
rect 707 705 819 717
rect 707 653 735 705
rect 787 653 819 705
rect 707 639 819 653
rect 986 798 1073 828
rect 986 746 1003 798
rect 1055 746 1073 798
rect 986 734 1073 746
rect 986 682 1003 734
rect 1055 682 1073 734
rect 986 652 1073 682
rect 1168 599 1202 844
rect 1059 598 1202 599
rect 479 555 1202 598
rect 1059 551 1202 555
rect -981 20 -889 28
rect -1108 -531 -1013 -54
rect -955 -318 -913 20
rect -881 -67 -816 -60
rect -881 -119 -874 -67
rect -822 -119 -816 -67
rect -881 -131 -816 -119
rect -881 -183 -874 -131
rect -822 -183 -816 -131
rect -881 -195 -816 -183
rect -881 -247 -874 -195
rect -822 -247 -816 -195
rect -881 -256 -816 -247
rect -685 -408 -580 54
rect -191 51 231 152
rect 10 13 122 51
rect -475 6 122 13
rect -523 -21 122 6
rect 325 -19 1114 16
rect -523 -317 -484 -21
rect -402 -255 -136 -59
rect -720 -413 -551 -408
rect -720 -465 -694 -413
rect -642 -465 -630 -413
rect -578 -465 -551 -413
rect -720 -469 -551 -465
rect -341 -531 -206 -255
rect -87 -317 -48 -21
rect 10 -257 122 -21
rect 244 -112 326 -78
rect 244 -164 257 -112
rect 309 -164 326 -112
rect 244 -176 326 -164
rect 244 -228 257 -176
rect 309 -228 326 -176
rect 244 -262 326 -228
rect 402 -92 484 -57
rect 402 -144 415 -92
rect 467 -144 484 -92
rect 402 -156 484 -144
rect 402 -208 415 -156
rect 467 -208 484 -156
rect 402 -241 484 -208
rect 563 -110 645 -76
rect 563 -162 576 -110
rect 628 -162 645 -110
rect 563 -174 645 -162
rect 563 -226 576 -174
rect 628 -226 645 -174
rect 563 -260 645 -226
rect 719 -92 801 -56
rect 719 -144 732 -92
rect 784 -144 801 -92
rect 719 -156 801 -144
rect 719 -208 732 -156
rect 784 -208 801 -156
rect 719 -240 801 -208
rect 879 -109 961 -74
rect 879 -161 894 -109
rect 946 -161 961 -109
rect 879 -173 961 -161
rect 879 -225 894 -173
rect 946 -225 961 -173
rect 879 -258 961 -225
rect 1028 -109 1114 -19
rect 1028 -161 1045 -109
rect 1097 -161 1114 -109
rect 1028 -173 1114 -161
rect 1028 -225 1045 -173
rect 1097 -225 1114 -173
rect 1028 -302 1114 -225
rect 1159 -257 1197 551
rect 1373 502 1404 1181
rect 1510 502 1553 1400
rect 1373 461 1553 502
rect 1911 489 1975 1505
rect 2534 1495 2683 1508
rect 1716 487 1975 489
rect 1716 435 1755 487
rect 1807 435 1819 487
rect 1871 435 1883 487
rect 1935 435 1975 487
rect 1716 434 1975 435
rect 2111 1402 2683 1445
rect 2111 1222 2147 1402
rect 2327 1222 2683 1402
rect 2111 1091 2683 1222
rect 1693 174 1726 175
rect 1583 122 1599 174
rect 1651 122 1663 174
rect 1715 122 1732 174
rect 1458 59 1529 78
rect 1458 15 1467 59
rect 1231 7 1467 15
rect 1519 7 1529 59
rect 1231 -5 1529 7
rect 1231 -15 1467 -5
rect 1458 -57 1467 -15
rect 1519 -57 1529 -5
rect 1458 -69 1529 -57
rect 1312 -107 1394 -72
rect 1312 -159 1327 -107
rect 1379 -159 1394 -107
rect 1312 -171 1394 -159
rect 1312 -223 1327 -171
rect 1379 -223 1394 -171
rect 1312 -256 1394 -223
rect 1458 -121 1467 -69
rect 1519 -121 1529 -69
rect 1458 -123 1529 -121
rect 1458 -133 1616 -123
rect 1458 -185 1467 -133
rect 1519 -185 1616 -133
rect 1458 -186 1616 -185
rect 1458 -197 1529 -186
rect 1458 -249 1467 -197
rect 1519 -249 1529 -197
rect 1458 -261 1529 -249
rect 1458 -302 1467 -261
rect 320 -313 1467 -302
rect 1519 -313 1529 -261
rect 1693 -308 1726 122
rect 320 -332 1529 -313
rect 1790 -367 1841 -54
rect 2111 -213 2363 1091
rect 2453 1002 2683 1026
rect 2453 694 2550 1002
rect 2666 694 2683 1002
rect 2453 588 2683 694
rect 2453 408 2478 588
rect 2658 408 2683 588
rect 2453 98 2683 408
rect 2453 -82 2478 98
rect 2658 -82 2683 98
rect 2453 -122 2683 -82
rect 2111 -283 2699 -213
rect 1790 -437 2589 -367
rect -4434 -701 -4382 -667
rect -4348 -701 -4296 -667
rect -4434 -739 -4296 -701
rect -4434 -773 -4382 -739
rect -4348 -773 -4296 -739
rect -4434 -811 -4296 -773
rect -4434 -845 -4382 -811
rect -4348 -845 -4296 -811
rect -4434 -883 -4296 -845
rect -4434 -917 -4382 -883
rect -4348 -917 -4296 -883
rect -4434 -955 -4296 -917
rect -4434 -989 -4382 -955
rect -4348 -989 -4296 -955
rect -4434 -1027 -4296 -989
rect -4434 -1061 -4382 -1027
rect -4348 -1061 -4296 -1027
rect -4434 -1099 -4296 -1061
rect -4434 -1133 -4382 -1099
rect -4348 -1133 -4296 -1099
rect -4434 -1171 -4296 -1133
rect -4434 -1205 -4382 -1171
rect -4348 -1205 -4296 -1171
rect -4434 -1243 -4296 -1205
rect -4434 -1277 -4382 -1243
rect -4348 -1277 -4296 -1243
rect -4434 -1315 -4296 -1277
rect -4434 -1349 -4382 -1315
rect -4348 -1349 -4296 -1315
rect -4434 -1387 -4296 -1349
rect -4434 -1421 -4382 -1387
rect -4348 -1421 -4296 -1387
rect -4434 -1459 -4296 -1421
rect -4434 -1493 -4382 -1459
rect -4348 -1493 -4296 -1459
rect -4434 -1531 -4296 -1493
rect -4434 -1565 -4382 -1531
rect -4348 -1565 -4296 -1531
rect -4434 -1603 -4296 -1565
rect -4434 -1637 -4382 -1603
rect -4348 -1637 -4296 -1603
rect -4434 -1675 -4296 -1637
rect -4434 -1709 -4382 -1675
rect -4348 -1709 -4296 -1675
rect -4434 -1747 -4296 -1709
rect -4434 -1781 -4382 -1747
rect -4348 -1781 -4296 -1747
rect -4434 -1819 -4296 -1781
rect -4434 -1853 -4382 -1819
rect -4348 -1853 -4296 -1819
rect -4434 -1891 -4296 -1853
rect -4434 -1925 -4382 -1891
rect -4348 -1925 -4296 -1891
rect -4434 -1963 -4296 -1925
rect -4434 -1997 -4382 -1963
rect -4348 -1997 -4296 -1963
rect -4434 -2055 -4296 -1997
rect -4196 -688 -3825 -621
rect -3707 -574 2271 -531
rect -3707 -626 -3657 -574
rect -3605 -626 -3593 -574
rect -3541 -626 -3529 -574
rect -3477 -583 -3465 -574
rect -3413 -583 -3401 -574
rect -3349 -583 -3337 -574
rect -3285 -583 -3273 -574
rect -3221 -583 -3209 -574
rect -3157 -583 -3145 -574
rect -3474 -617 -3465 -583
rect -3402 -617 -3401 -583
rect -3221 -617 -3220 -583
rect -3157 -617 -3148 -583
rect -3477 -626 -3465 -617
rect -3413 -626 -3401 -617
rect -3349 -626 -3337 -617
rect -3285 -626 -3273 -617
rect -3221 -626 -3209 -617
rect -3157 -626 -3145 -617
rect -3093 -626 -3081 -574
rect -3029 -626 -3017 -574
rect -2965 -626 -2953 -574
rect -2901 -583 -2889 -574
rect -2837 -583 -2825 -574
rect -2773 -583 -2761 -574
rect -2709 -583 -2697 -574
rect -2645 -583 -2633 -574
rect -2581 -583 -2569 -574
rect -2898 -617 -2889 -583
rect -2826 -617 -2825 -583
rect -2645 -617 -2644 -583
rect -2581 -617 -2572 -583
rect -2901 -626 -2889 -617
rect -2837 -626 -2825 -617
rect -2773 -626 -2761 -617
rect -2709 -626 -2697 -617
rect -2645 -626 -2633 -617
rect -2581 -626 -2569 -617
rect -2517 -626 -2505 -574
rect -2453 -626 -2441 -574
rect -2389 -626 -2377 -574
rect -2325 -583 -2313 -574
rect -2261 -583 -2249 -574
rect -2197 -583 -2185 -574
rect -2133 -583 -2121 -574
rect -2069 -583 -2057 -574
rect -2005 -583 -1993 -574
rect -2322 -617 -2313 -583
rect -2250 -617 -2249 -583
rect -2069 -617 -2068 -583
rect -2005 -617 -1996 -583
rect -2325 -626 -2313 -617
rect -2261 -626 -2249 -617
rect -2197 -626 -2185 -617
rect -2133 -626 -2121 -617
rect -2069 -626 -2057 -617
rect -2005 -626 -1993 -617
rect -1941 -626 -1929 -574
rect -1877 -626 -1865 -574
rect -1813 -626 -1801 -574
rect -1749 -583 -1737 -574
rect -1685 -583 -1673 -574
rect -1621 -583 -1609 -574
rect -1557 -583 -1545 -574
rect -1493 -583 -1481 -574
rect -1429 -583 -1417 -574
rect -1746 -617 -1737 -583
rect -1674 -617 -1673 -583
rect -1493 -617 -1492 -583
rect -1429 -617 -1420 -583
rect -1749 -626 -1737 -617
rect -1685 -626 -1673 -617
rect -1621 -626 -1609 -617
rect -1557 -626 -1545 -617
rect -1493 -626 -1481 -617
rect -1429 -626 -1417 -617
rect -1365 -626 -1353 -574
rect -1301 -626 -1289 -574
rect -1237 -626 -1225 -574
rect -1173 -583 -1161 -574
rect -1109 -583 -1097 -574
rect -1045 -583 -1033 -574
rect -981 -583 -969 -574
rect -917 -583 -905 -574
rect -853 -583 -841 -574
rect -1170 -617 -1161 -583
rect -1098 -617 -1097 -583
rect -917 -617 -916 -583
rect -853 -617 -844 -583
rect -1173 -626 -1161 -617
rect -1109 -626 -1097 -617
rect -1045 -626 -1033 -617
rect -981 -626 -969 -617
rect -917 -626 -905 -617
rect -853 -626 -841 -617
rect -789 -626 -777 -574
rect -725 -626 -713 -574
rect -661 -626 -649 -574
rect -597 -583 -585 -574
rect -533 -583 -521 -574
rect -469 -583 -457 -574
rect -405 -583 -393 -574
rect -341 -583 -329 -574
rect -277 -583 -265 -574
rect -594 -617 -585 -583
rect -522 -617 -521 -583
rect -341 -617 -340 -583
rect -277 -617 -268 -583
rect -597 -626 -585 -617
rect -533 -626 -521 -617
rect -469 -626 -457 -617
rect -405 -626 -393 -617
rect -341 -626 -329 -617
rect -277 -626 -265 -617
rect -213 -626 -201 -574
rect -149 -626 -137 -574
rect -85 -626 -73 -574
rect -21 -583 -9 -574
rect 43 -583 55 -574
rect 107 -583 119 -574
rect 171 -583 183 -574
rect 235 -583 247 -574
rect 299 -583 311 -574
rect -18 -617 -9 -583
rect 54 -617 55 -583
rect 235 -617 236 -583
rect 299 -617 308 -583
rect -21 -626 -9 -617
rect 43 -626 55 -617
rect 107 -626 119 -617
rect 171 -626 183 -617
rect 235 -626 247 -617
rect 299 -626 311 -617
rect 363 -626 375 -574
rect 427 -626 439 -574
rect 491 -626 503 -574
rect 555 -583 567 -574
rect 619 -583 631 -574
rect 683 -583 695 -574
rect 747 -583 759 -574
rect 811 -583 823 -574
rect 875 -583 887 -574
rect 558 -617 567 -583
rect 630 -617 631 -583
rect 811 -617 812 -583
rect 875 -617 884 -583
rect 555 -626 567 -617
rect 619 -626 631 -617
rect 683 -626 695 -617
rect 747 -626 759 -617
rect 811 -626 823 -617
rect 875 -626 887 -617
rect 939 -626 951 -574
rect 1003 -626 1015 -574
rect 1067 -626 1079 -574
rect 1131 -583 1143 -574
rect 1195 -583 1207 -574
rect 1259 -583 1271 -574
rect 1323 -583 1335 -574
rect 1387 -583 1399 -574
rect 1451 -583 1463 -574
rect 1134 -617 1143 -583
rect 1206 -617 1207 -583
rect 1387 -617 1388 -583
rect 1451 -617 1460 -583
rect 1131 -626 1143 -617
rect 1195 -626 1207 -617
rect 1259 -626 1271 -617
rect 1323 -626 1335 -617
rect 1387 -626 1399 -617
rect 1451 -626 1463 -617
rect 1515 -626 1527 -574
rect 1579 -626 1591 -574
rect 1643 -626 1655 -574
rect 1707 -583 1719 -574
rect 1771 -583 1783 -574
rect 1835 -583 1847 -574
rect 1899 -583 1911 -574
rect 1963 -583 1975 -574
rect 2027 -583 2039 -574
rect 1710 -617 1719 -583
rect 1782 -617 1783 -583
rect 1963 -617 1964 -583
rect 2027 -617 2036 -583
rect 1707 -626 1719 -617
rect 1771 -626 1783 -617
rect 1835 -626 1847 -617
rect 1899 -626 1911 -617
rect 1963 -626 1975 -617
rect 2027 -626 2039 -617
rect 2091 -626 2103 -574
rect 2155 -626 2167 -574
rect 2219 -626 2271 -574
rect -3707 -660 2271 -626
rect -4196 -756 -4129 -688
rect -4196 -823 2475 -756
rect -4196 -1125 -4129 -823
rect -4072 -884 -3944 -878
rect -4072 -936 -4066 -884
rect -4014 -936 -4002 -884
rect -3950 -936 -3944 -884
rect -4072 -942 -3944 -936
rect -3756 -884 -3628 -878
rect -3756 -936 -3750 -884
rect -3698 -936 -3686 -884
rect -3634 -936 -3628 -884
rect -3756 -942 -3628 -936
rect -3440 -884 -3312 -878
rect -3440 -936 -3434 -884
rect -3382 -936 -3370 -884
rect -3318 -936 -3312 -884
rect -3440 -942 -3312 -936
rect -3124 -884 -2996 -878
rect -3124 -936 -3118 -884
rect -3066 -936 -3054 -884
rect -3002 -936 -2996 -884
rect -3124 -942 -2996 -936
rect -2808 -884 -2680 -878
rect -2808 -936 -2802 -884
rect -2750 -936 -2738 -884
rect -2686 -936 -2680 -884
rect -2808 -942 -2680 -936
rect -2492 -884 -2364 -878
rect -2492 -936 -2486 -884
rect -2434 -936 -2422 -884
rect -2370 -936 -2364 -884
rect -2492 -942 -2364 -936
rect -2176 -884 -2048 -878
rect -2176 -936 -2170 -884
rect -2118 -936 -2106 -884
rect -2054 -936 -2048 -884
rect -2176 -942 -2048 -936
rect -1860 -884 -1732 -878
rect -1860 -936 -1854 -884
rect -1802 -936 -1790 -884
rect -1738 -936 -1732 -884
rect -1860 -942 -1732 -936
rect -1544 -884 -1416 -878
rect -1544 -936 -1538 -884
rect -1486 -936 -1474 -884
rect -1422 -936 -1416 -884
rect -1544 -942 -1416 -936
rect -1228 -884 -1100 -878
rect -1228 -936 -1222 -884
rect -1170 -936 -1158 -884
rect -1106 -936 -1100 -884
rect -1228 -942 -1100 -936
rect -912 -884 -784 -878
rect -912 -936 -906 -884
rect -854 -936 -842 -884
rect -790 -936 -784 -884
rect -912 -942 -784 -936
rect -596 -884 -468 -878
rect -596 -936 -590 -884
rect -538 -936 -526 -884
rect -474 -936 -468 -884
rect -596 -942 -468 -936
rect -280 -884 -152 -878
rect -280 -936 -274 -884
rect -222 -936 -210 -884
rect -158 -936 -152 -884
rect -280 -942 -152 -936
rect 36 -884 164 -878
rect 36 -936 42 -884
rect 94 -936 106 -884
rect 158 -936 164 -884
rect 36 -942 164 -936
rect 352 -884 480 -878
rect 352 -936 358 -884
rect 410 -936 422 -884
rect 474 -936 480 -884
rect 352 -942 480 -936
rect 668 -884 796 -878
rect 668 -936 674 -884
rect 726 -936 738 -884
rect 790 -936 796 -884
rect 668 -942 796 -936
rect 984 -884 1112 -878
rect 984 -936 990 -884
rect 1042 -936 1054 -884
rect 1106 -936 1112 -884
rect 984 -942 1112 -936
rect 1300 -884 1428 -878
rect 1300 -936 1306 -884
rect 1358 -936 1370 -884
rect 1422 -936 1428 -884
rect 1300 -942 1428 -936
rect 1616 -884 1744 -878
rect 1616 -936 1622 -884
rect 1674 -936 1686 -884
rect 1738 -936 1744 -884
rect 1616 -942 1744 -936
rect 1932 -884 2060 -878
rect 1932 -936 1938 -884
rect 1990 -936 2002 -884
rect 2054 -936 2060 -884
rect 1932 -942 2060 -936
rect 2248 -884 2376 -878
rect 2248 -936 2254 -884
rect 2306 -936 2318 -884
rect 2370 -936 2376 -884
rect 2248 -942 2376 -936
rect -3914 -1009 -3786 -1003
rect -3914 -1061 -3908 -1009
rect -3856 -1061 -3844 -1009
rect -3792 -1061 -3786 -1009
rect -3914 -1067 -3786 -1061
rect -3598 -1009 -3470 -1003
rect -3598 -1061 -3592 -1009
rect -3540 -1061 -3528 -1009
rect -3476 -1061 -3470 -1009
rect -3598 -1067 -3470 -1061
rect -3282 -1009 -3154 -1003
rect -3282 -1061 -3276 -1009
rect -3224 -1061 -3212 -1009
rect -3160 -1061 -3154 -1009
rect -3282 -1067 -3154 -1061
rect -2966 -1009 -2838 -1003
rect -2966 -1061 -2960 -1009
rect -2908 -1061 -2896 -1009
rect -2844 -1061 -2838 -1009
rect -2966 -1067 -2838 -1061
rect -2650 -1009 -2522 -1003
rect -2650 -1061 -2644 -1009
rect -2592 -1061 -2580 -1009
rect -2528 -1061 -2522 -1009
rect -2650 -1067 -2522 -1061
rect -2334 -1009 -2206 -1003
rect -2334 -1061 -2328 -1009
rect -2276 -1061 -2264 -1009
rect -2212 -1061 -2206 -1009
rect -2334 -1067 -2206 -1061
rect -2018 -1009 -1890 -1003
rect -2018 -1061 -2012 -1009
rect -1960 -1061 -1948 -1009
rect -1896 -1061 -1890 -1009
rect -2018 -1067 -1890 -1061
rect -1702 -1009 -1574 -1003
rect -1702 -1061 -1696 -1009
rect -1644 -1061 -1632 -1009
rect -1580 -1061 -1574 -1009
rect -1702 -1067 -1574 -1061
rect -1386 -1009 -1258 -1003
rect -1386 -1061 -1380 -1009
rect -1328 -1061 -1316 -1009
rect -1264 -1061 -1258 -1009
rect -1386 -1067 -1258 -1061
rect -1070 -1009 -942 -1003
rect -1070 -1061 -1064 -1009
rect -1012 -1061 -1000 -1009
rect -948 -1061 -942 -1009
rect -1070 -1067 -942 -1061
rect -754 -1009 -626 -1003
rect -754 -1061 -748 -1009
rect -696 -1061 -684 -1009
rect -632 -1061 -626 -1009
rect -754 -1067 -626 -1061
rect -438 -1009 -310 -1003
rect -438 -1061 -432 -1009
rect -380 -1061 -368 -1009
rect -316 -1061 -310 -1009
rect -438 -1067 -310 -1061
rect -122 -1009 6 -1003
rect -122 -1061 -116 -1009
rect -64 -1061 -52 -1009
rect 0 -1061 6 -1009
rect -122 -1067 6 -1061
rect 194 -1009 322 -1003
rect 194 -1061 200 -1009
rect 252 -1061 264 -1009
rect 316 -1061 322 -1009
rect 194 -1067 322 -1061
rect 510 -1009 638 -1003
rect 510 -1061 516 -1009
rect 568 -1061 580 -1009
rect 632 -1061 638 -1009
rect 510 -1067 638 -1061
rect 826 -1009 954 -1003
rect 826 -1061 832 -1009
rect 884 -1061 896 -1009
rect 948 -1061 954 -1009
rect 826 -1067 954 -1061
rect 1142 -1009 1270 -1003
rect 1142 -1061 1148 -1009
rect 1200 -1061 1212 -1009
rect 1264 -1061 1270 -1009
rect 1142 -1067 1270 -1061
rect 1458 -1009 1586 -1003
rect 1458 -1061 1464 -1009
rect 1516 -1061 1528 -1009
rect 1580 -1061 1586 -1009
rect 1458 -1067 1586 -1061
rect 1774 -1009 1902 -1003
rect 1774 -1061 1780 -1009
rect 1832 -1061 1844 -1009
rect 1896 -1061 1902 -1009
rect 1774 -1067 1902 -1061
rect 2090 -1009 2218 -1003
rect 2090 -1061 2096 -1009
rect 2148 -1061 2160 -1009
rect 2212 -1061 2218 -1009
rect 2090 -1067 2218 -1061
rect 2408 -1125 2475 -823
rect -4196 -1240 2475 -1125
rect -4196 -1546 -4129 -1240
rect -4072 -1302 -3944 -1296
rect -4072 -1354 -4066 -1302
rect -4014 -1354 -4002 -1302
rect -3950 -1354 -3944 -1302
rect -4072 -1360 -3944 -1354
rect -3756 -1302 -3628 -1296
rect -3756 -1354 -3750 -1302
rect -3698 -1354 -3686 -1302
rect -3634 -1354 -3628 -1302
rect -3756 -1360 -3628 -1354
rect -3440 -1302 -3312 -1296
rect -3440 -1354 -3434 -1302
rect -3382 -1354 -3370 -1302
rect -3318 -1354 -3312 -1302
rect -3440 -1360 -3312 -1354
rect -3124 -1302 -2996 -1296
rect -3124 -1354 -3118 -1302
rect -3066 -1354 -3054 -1302
rect -3002 -1354 -2996 -1302
rect -3124 -1360 -2996 -1354
rect -2808 -1302 -2680 -1296
rect -2808 -1354 -2802 -1302
rect -2750 -1354 -2738 -1302
rect -2686 -1354 -2680 -1302
rect -2808 -1360 -2680 -1354
rect -2492 -1302 -2364 -1296
rect -2492 -1354 -2486 -1302
rect -2434 -1354 -2422 -1302
rect -2370 -1354 -2364 -1302
rect -2492 -1360 -2364 -1354
rect -2176 -1302 -2048 -1296
rect -2176 -1354 -2170 -1302
rect -2118 -1354 -2106 -1302
rect -2054 -1354 -2048 -1302
rect -2176 -1360 -2048 -1354
rect -1860 -1302 -1732 -1296
rect -1860 -1354 -1854 -1302
rect -1802 -1354 -1790 -1302
rect -1738 -1354 -1732 -1302
rect -1860 -1360 -1732 -1354
rect -1544 -1302 -1416 -1296
rect -1544 -1354 -1538 -1302
rect -1486 -1354 -1474 -1302
rect -1422 -1354 -1416 -1302
rect -1544 -1360 -1416 -1354
rect -1228 -1302 -1100 -1296
rect -1228 -1354 -1222 -1302
rect -1170 -1354 -1158 -1302
rect -1106 -1354 -1100 -1302
rect -1228 -1360 -1100 -1354
rect -912 -1302 -784 -1296
rect -912 -1354 -906 -1302
rect -854 -1354 -842 -1302
rect -790 -1354 -784 -1302
rect -912 -1360 -784 -1354
rect -596 -1302 -468 -1296
rect -596 -1354 -590 -1302
rect -538 -1354 -526 -1302
rect -474 -1354 -468 -1302
rect -596 -1360 -468 -1354
rect -280 -1302 -152 -1296
rect -280 -1354 -274 -1302
rect -222 -1354 -210 -1302
rect -158 -1354 -152 -1302
rect -280 -1360 -152 -1354
rect 36 -1302 164 -1296
rect 36 -1354 42 -1302
rect 94 -1354 106 -1302
rect 158 -1354 164 -1302
rect 36 -1360 164 -1354
rect 352 -1302 480 -1296
rect 352 -1354 358 -1302
rect 410 -1354 422 -1302
rect 474 -1354 480 -1302
rect 352 -1360 480 -1354
rect 668 -1302 796 -1296
rect 668 -1354 674 -1302
rect 726 -1354 738 -1302
rect 790 -1354 796 -1302
rect 668 -1360 796 -1354
rect 984 -1302 1112 -1296
rect 984 -1354 990 -1302
rect 1042 -1354 1054 -1302
rect 1106 -1354 1112 -1302
rect 984 -1360 1112 -1354
rect 1300 -1302 1428 -1296
rect 1300 -1354 1306 -1302
rect 1358 -1354 1370 -1302
rect 1422 -1354 1428 -1302
rect 1300 -1360 1428 -1354
rect 1616 -1302 1744 -1296
rect 1616 -1354 1622 -1302
rect 1674 -1354 1686 -1302
rect 1738 -1354 1744 -1302
rect 1616 -1360 1744 -1354
rect 1932 -1302 2060 -1296
rect 1932 -1354 1938 -1302
rect 1990 -1354 2002 -1302
rect 2054 -1354 2060 -1302
rect 1932 -1360 2060 -1354
rect 2248 -1302 2376 -1296
rect 2248 -1354 2254 -1302
rect 2306 -1354 2318 -1302
rect 2370 -1354 2376 -1302
rect 2248 -1360 2376 -1354
rect -3914 -1427 -3786 -1421
rect -3914 -1479 -3908 -1427
rect -3856 -1479 -3844 -1427
rect -3792 -1479 -3786 -1427
rect -3914 -1485 -3786 -1479
rect -3598 -1427 -3470 -1421
rect -3598 -1479 -3592 -1427
rect -3540 -1479 -3528 -1427
rect -3476 -1479 -3470 -1427
rect -3598 -1485 -3470 -1479
rect -3282 -1427 -3154 -1421
rect -3282 -1479 -3276 -1427
rect -3224 -1479 -3212 -1427
rect -3160 -1479 -3154 -1427
rect -3282 -1485 -3154 -1479
rect -2966 -1427 -2838 -1421
rect -2966 -1479 -2960 -1427
rect -2908 -1479 -2896 -1427
rect -2844 -1479 -2838 -1427
rect -2966 -1485 -2838 -1479
rect -2650 -1427 -2522 -1421
rect -2650 -1479 -2644 -1427
rect -2592 -1479 -2580 -1427
rect -2528 -1479 -2522 -1427
rect -2650 -1485 -2522 -1479
rect -2334 -1427 -2206 -1421
rect -2334 -1479 -2328 -1427
rect -2276 -1479 -2264 -1427
rect -2212 -1479 -2206 -1427
rect -2334 -1485 -2206 -1479
rect -2018 -1427 -1890 -1421
rect -2018 -1479 -2012 -1427
rect -1960 -1479 -1948 -1427
rect -1896 -1479 -1890 -1427
rect -2018 -1485 -1890 -1479
rect -1702 -1427 -1574 -1421
rect -1702 -1479 -1696 -1427
rect -1644 -1479 -1632 -1427
rect -1580 -1479 -1574 -1427
rect -1702 -1485 -1574 -1479
rect -1386 -1427 -1258 -1421
rect -1386 -1479 -1380 -1427
rect -1328 -1479 -1316 -1427
rect -1264 -1479 -1258 -1427
rect -1386 -1485 -1258 -1479
rect -1070 -1427 -942 -1421
rect -1070 -1479 -1064 -1427
rect -1012 -1479 -1000 -1427
rect -948 -1479 -942 -1427
rect -1070 -1485 -942 -1479
rect -754 -1427 -626 -1421
rect -754 -1479 -748 -1427
rect -696 -1479 -684 -1427
rect -632 -1479 -626 -1427
rect -754 -1485 -626 -1479
rect -438 -1427 -310 -1421
rect -438 -1479 -432 -1427
rect -380 -1479 -368 -1427
rect -316 -1479 -310 -1427
rect -438 -1485 -310 -1479
rect -122 -1427 6 -1421
rect -122 -1479 -116 -1427
rect -64 -1479 -52 -1427
rect 0 -1479 6 -1427
rect -122 -1485 6 -1479
rect 194 -1427 322 -1421
rect 194 -1479 200 -1427
rect 252 -1479 264 -1427
rect 316 -1479 322 -1427
rect 194 -1485 322 -1479
rect 510 -1427 638 -1421
rect 510 -1479 516 -1427
rect 568 -1479 580 -1427
rect 632 -1479 638 -1427
rect 510 -1485 638 -1479
rect 826 -1427 954 -1421
rect 826 -1479 832 -1427
rect 884 -1479 896 -1427
rect 948 -1479 954 -1427
rect 826 -1485 954 -1479
rect 1142 -1427 1270 -1421
rect 1142 -1479 1148 -1427
rect 1200 -1479 1212 -1427
rect 1264 -1479 1270 -1427
rect 1142 -1485 1270 -1479
rect 1458 -1427 1586 -1421
rect 1458 -1479 1464 -1427
rect 1516 -1479 1528 -1427
rect 1580 -1479 1586 -1427
rect 1458 -1485 1586 -1479
rect 1774 -1427 1902 -1421
rect 1774 -1479 1780 -1427
rect 1832 -1479 1844 -1427
rect 1896 -1479 1902 -1427
rect 1774 -1485 1902 -1479
rect 2090 -1427 2218 -1421
rect 2090 -1479 2096 -1427
rect 2148 -1479 2160 -1427
rect 2212 -1479 2218 -1427
rect 2090 -1485 2218 -1479
rect 2408 -1546 2475 -1240
rect -4196 -1661 2475 -1546
rect -4196 -1956 -4129 -1661
rect -4072 -1720 -3944 -1714
rect -4072 -1772 -4066 -1720
rect -4014 -1772 -4002 -1720
rect -3950 -1772 -3944 -1720
rect -4072 -1778 -3944 -1772
rect -3756 -1720 -3628 -1714
rect -3756 -1772 -3750 -1720
rect -3698 -1772 -3686 -1720
rect -3634 -1772 -3628 -1720
rect -3756 -1778 -3628 -1772
rect -3440 -1720 -3312 -1714
rect -3440 -1772 -3434 -1720
rect -3382 -1772 -3370 -1720
rect -3318 -1772 -3312 -1720
rect -3440 -1778 -3312 -1772
rect -3124 -1720 -2996 -1714
rect -3124 -1772 -3118 -1720
rect -3066 -1772 -3054 -1720
rect -3002 -1772 -2996 -1720
rect -3124 -1778 -2996 -1772
rect -2808 -1720 -2680 -1714
rect -2808 -1772 -2802 -1720
rect -2750 -1772 -2738 -1720
rect -2686 -1772 -2680 -1720
rect -2808 -1778 -2680 -1772
rect -2492 -1720 -2364 -1714
rect -2492 -1772 -2486 -1720
rect -2434 -1772 -2422 -1720
rect -2370 -1772 -2364 -1720
rect -2492 -1778 -2364 -1772
rect -2176 -1720 -2048 -1714
rect -2176 -1772 -2170 -1720
rect -2118 -1772 -2106 -1720
rect -2054 -1772 -2048 -1720
rect -2176 -1778 -2048 -1772
rect -1860 -1720 -1732 -1714
rect -1860 -1772 -1854 -1720
rect -1802 -1772 -1790 -1720
rect -1738 -1772 -1732 -1720
rect -1860 -1778 -1732 -1772
rect -1544 -1720 -1416 -1714
rect -1544 -1772 -1538 -1720
rect -1486 -1772 -1474 -1720
rect -1422 -1772 -1416 -1720
rect -1544 -1778 -1416 -1772
rect -1228 -1720 -1100 -1714
rect -1228 -1772 -1222 -1720
rect -1170 -1772 -1158 -1720
rect -1106 -1772 -1100 -1720
rect -1228 -1778 -1100 -1772
rect -912 -1720 -784 -1714
rect -912 -1772 -906 -1720
rect -854 -1772 -842 -1720
rect -790 -1772 -784 -1720
rect -912 -1778 -784 -1772
rect -596 -1720 -468 -1714
rect -596 -1772 -590 -1720
rect -538 -1772 -526 -1720
rect -474 -1772 -468 -1720
rect -596 -1778 -468 -1772
rect -280 -1720 -152 -1714
rect -280 -1772 -274 -1720
rect -222 -1772 -210 -1720
rect -158 -1772 -152 -1720
rect -280 -1778 -152 -1772
rect 36 -1720 164 -1714
rect 36 -1772 42 -1720
rect 94 -1772 106 -1720
rect 158 -1772 164 -1720
rect 36 -1778 164 -1772
rect 352 -1720 480 -1714
rect 352 -1772 358 -1720
rect 410 -1772 422 -1720
rect 474 -1772 480 -1720
rect 352 -1778 480 -1772
rect 668 -1720 796 -1714
rect 668 -1772 674 -1720
rect 726 -1772 738 -1720
rect 790 -1772 796 -1720
rect 668 -1778 796 -1772
rect 984 -1720 1112 -1714
rect 984 -1772 990 -1720
rect 1042 -1772 1054 -1720
rect 1106 -1772 1112 -1720
rect 984 -1778 1112 -1772
rect 1300 -1720 1428 -1714
rect 1300 -1772 1306 -1720
rect 1358 -1772 1370 -1720
rect 1422 -1772 1428 -1720
rect 1300 -1778 1428 -1772
rect 1616 -1720 1744 -1714
rect 1616 -1772 1622 -1720
rect 1674 -1772 1686 -1720
rect 1738 -1772 1744 -1720
rect 1616 -1778 1744 -1772
rect 1932 -1720 2060 -1714
rect 1932 -1772 1938 -1720
rect 1990 -1772 2002 -1720
rect 2054 -1772 2060 -1720
rect 1932 -1778 2060 -1772
rect 2248 -1720 2376 -1714
rect 2248 -1772 2254 -1720
rect 2306 -1772 2318 -1720
rect 2370 -1772 2376 -1720
rect 2248 -1778 2376 -1772
rect -3914 -1845 -3786 -1839
rect -3914 -1897 -3908 -1845
rect -3856 -1897 -3844 -1845
rect -3792 -1897 -3786 -1845
rect -3914 -1903 -3786 -1897
rect -3598 -1845 -3470 -1839
rect -3598 -1897 -3592 -1845
rect -3540 -1897 -3528 -1845
rect -3476 -1897 -3470 -1845
rect -3598 -1903 -3470 -1897
rect -3282 -1845 -3154 -1839
rect -3282 -1897 -3276 -1845
rect -3224 -1897 -3212 -1845
rect -3160 -1897 -3154 -1845
rect -3282 -1903 -3154 -1897
rect -2966 -1845 -2838 -1839
rect -2966 -1897 -2960 -1845
rect -2908 -1897 -2896 -1845
rect -2844 -1897 -2838 -1845
rect -2966 -1903 -2838 -1897
rect -2650 -1845 -2522 -1839
rect -2650 -1897 -2644 -1845
rect -2592 -1897 -2580 -1845
rect -2528 -1897 -2522 -1845
rect -2650 -1903 -2522 -1897
rect -2334 -1845 -2206 -1839
rect -2334 -1897 -2328 -1845
rect -2276 -1897 -2264 -1845
rect -2212 -1897 -2206 -1845
rect -2334 -1903 -2206 -1897
rect -2018 -1845 -1890 -1839
rect -2018 -1897 -2012 -1845
rect -1960 -1897 -1948 -1845
rect -1896 -1897 -1890 -1845
rect -2018 -1903 -1890 -1897
rect -1702 -1845 -1574 -1839
rect -1702 -1897 -1696 -1845
rect -1644 -1897 -1632 -1845
rect -1580 -1897 -1574 -1845
rect -1702 -1903 -1574 -1897
rect -1386 -1845 -1258 -1839
rect -1386 -1897 -1380 -1845
rect -1328 -1897 -1316 -1845
rect -1264 -1897 -1258 -1845
rect -1386 -1903 -1258 -1897
rect -1070 -1845 -942 -1839
rect -1070 -1897 -1064 -1845
rect -1012 -1897 -1000 -1845
rect -948 -1897 -942 -1845
rect -1070 -1903 -942 -1897
rect -754 -1845 -626 -1839
rect -754 -1897 -748 -1845
rect -696 -1897 -684 -1845
rect -632 -1897 -626 -1845
rect -754 -1903 -626 -1897
rect -438 -1845 -310 -1839
rect -438 -1897 -432 -1845
rect -380 -1897 -368 -1845
rect -316 -1897 -310 -1845
rect -438 -1903 -310 -1897
rect -122 -1845 6 -1839
rect -122 -1897 -116 -1845
rect -64 -1897 -52 -1845
rect 0 -1897 6 -1845
rect -122 -1903 6 -1897
rect 194 -1845 322 -1839
rect 194 -1897 200 -1845
rect 252 -1897 264 -1845
rect 316 -1897 322 -1845
rect 194 -1903 322 -1897
rect 510 -1845 638 -1839
rect 510 -1897 516 -1845
rect 568 -1897 580 -1845
rect 632 -1897 638 -1845
rect 510 -1903 638 -1897
rect 826 -1845 954 -1839
rect 826 -1897 832 -1845
rect 884 -1897 896 -1845
rect 948 -1897 954 -1845
rect 826 -1903 954 -1897
rect 1142 -1845 1270 -1839
rect 1142 -1897 1148 -1845
rect 1200 -1897 1212 -1845
rect 1264 -1897 1270 -1845
rect 1142 -1903 1270 -1897
rect 1458 -1845 1586 -1839
rect 1458 -1897 1464 -1845
rect 1516 -1897 1528 -1845
rect 1580 -1897 1586 -1845
rect 1458 -1903 1586 -1897
rect 1774 -1845 1902 -1839
rect 1774 -1897 1780 -1845
rect 1832 -1897 1844 -1845
rect 1896 -1897 1902 -1845
rect 1774 -1903 1902 -1897
rect 2090 -1845 2218 -1839
rect 2090 -1897 2096 -1845
rect 2148 -1897 2160 -1845
rect 2212 -1897 2218 -1845
rect 2090 -1903 2218 -1897
rect 2408 -1956 2475 -1661
rect -4196 -2023 2475 -1956
rect -4392 -2131 2353 -2099
rect -4392 -2439 -4380 -2131
rect -4136 -2167 2353 -2131
rect -4136 -2173 -3897 -2167
rect -4136 -2207 -4079 -2173
rect -4045 -2201 -3897 -2173
rect -3863 -2201 -3825 -2167
rect -3791 -2201 -3753 -2167
rect -3719 -2201 -3681 -2167
rect -3647 -2201 -3609 -2167
rect -3575 -2201 -3537 -2167
rect -3503 -2201 -3465 -2167
rect -3431 -2201 -3393 -2167
rect -3359 -2201 -3321 -2167
rect -3287 -2201 -3249 -2167
rect -3215 -2201 -3177 -2167
rect -3143 -2201 -3105 -2167
rect -3071 -2201 -3033 -2167
rect -2999 -2201 -2961 -2167
rect -2927 -2201 -2889 -2167
rect -2855 -2201 -2817 -2167
rect -2783 -2201 -2745 -2167
rect -2711 -2201 -2673 -2167
rect -2639 -2201 -2601 -2167
rect -2567 -2201 -2529 -2167
rect -2495 -2201 -2457 -2167
rect -2423 -2201 -2385 -2167
rect -2351 -2201 -2313 -2167
rect -2279 -2201 -2241 -2167
rect -2207 -2201 -2169 -2167
rect -2135 -2201 -2097 -2167
rect -2063 -2201 -2025 -2167
rect -1991 -2201 -1953 -2167
rect -1919 -2201 -1881 -2167
rect -1847 -2201 -1809 -2167
rect -1775 -2201 -1737 -2167
rect -1703 -2201 -1665 -2167
rect -1631 -2201 -1593 -2167
rect -1559 -2201 -1521 -2167
rect -1487 -2201 -1449 -2167
rect -1415 -2201 -1377 -2167
rect -1343 -2201 -1305 -2167
rect -1271 -2201 -1233 -2167
rect -1199 -2201 -1161 -2167
rect -1127 -2201 -1089 -2167
rect -1055 -2201 -1017 -2167
rect -983 -2201 -945 -2167
rect -911 -2201 -873 -2167
rect -839 -2201 -801 -2167
rect -767 -2201 -729 -2167
rect -695 -2201 -657 -2167
rect -623 -2201 -585 -2167
rect -551 -2201 -513 -2167
rect -479 -2201 -441 -2167
rect -407 -2201 -369 -2167
rect -335 -2201 -297 -2167
rect -263 -2201 -225 -2167
rect -191 -2201 -153 -2167
rect -119 -2201 -81 -2167
rect -47 -2201 -9 -2167
rect 25 -2201 63 -2167
rect 97 -2201 135 -2167
rect 169 -2201 207 -2167
rect 241 -2201 279 -2167
rect 313 -2201 351 -2167
rect 385 -2201 423 -2167
rect 457 -2201 495 -2167
rect 529 -2201 567 -2167
rect 601 -2201 639 -2167
rect 673 -2201 711 -2167
rect 745 -2201 783 -2167
rect 817 -2201 855 -2167
rect 889 -2201 927 -2167
rect 961 -2201 999 -2167
rect 1033 -2201 1071 -2167
rect 1105 -2201 1143 -2167
rect 1177 -2201 1215 -2167
rect 1249 -2201 1287 -2167
rect 1321 -2201 1359 -2167
rect 1393 -2201 1431 -2167
rect 1465 -2201 1503 -2167
rect 1537 -2201 1575 -2167
rect 1609 -2201 1647 -2167
rect 1681 -2201 1719 -2167
rect 1753 -2201 1791 -2167
rect 1825 -2201 1863 -2167
rect 1897 -2201 1935 -2167
rect 1969 -2201 2007 -2167
rect 2041 -2201 2079 -2167
rect 2113 -2201 2151 -2167
rect 2185 -2201 2223 -2167
rect 2257 -2201 2295 -2167
rect 2329 -2201 2353 -2167
rect -4045 -2207 2353 -2201
rect -4136 -2245 2353 -2207
rect -4136 -2279 -4079 -2245
rect -4045 -2255 2353 -2245
rect -4045 -2279 -3994 -2255
rect -4136 -2317 -3994 -2279
rect -4136 -2351 -4079 -2317
rect -4045 -2351 -3994 -2317
rect -4136 -2389 -3994 -2351
rect -4136 -2423 -4079 -2389
rect -4045 -2423 -3994 -2389
rect -4136 -2439 -3994 -2423
rect -4392 -2461 -3994 -2439
rect -4392 -2472 -4079 -2461
rect -4125 -2495 -4079 -2472
rect -4045 -2495 -3994 -2461
rect -4125 -2533 -3994 -2495
rect -4434 -2618 -4296 -2548
rect -4434 -2652 -4375 -2618
rect -4341 -2652 -4296 -2618
rect -4434 -2690 -4296 -2652
rect -4434 -2724 -4375 -2690
rect -4341 -2724 -4296 -2690
rect -4434 -2762 -4296 -2724
rect -4434 -2796 -4375 -2762
rect -4341 -2796 -4296 -2762
rect -4434 -2834 -4296 -2796
rect -4434 -2868 -4375 -2834
rect -4341 -2868 -4296 -2834
rect -4434 -2906 -4296 -2868
rect -4434 -2940 -4375 -2906
rect -4341 -2940 -4296 -2906
rect -4434 -2978 -4296 -2940
rect -4434 -3012 -4375 -2978
rect -4341 -3012 -4296 -2978
rect -4434 -3050 -4296 -3012
rect -4434 -3084 -4375 -3050
rect -4341 -3084 -4296 -3050
rect -4434 -3122 -4296 -3084
rect -4434 -3156 -4375 -3122
rect -4341 -3156 -4296 -3122
rect -4434 -3194 -4296 -3156
rect -4434 -3228 -4375 -3194
rect -4341 -3228 -4296 -3194
rect -4434 -3266 -4296 -3228
rect -4434 -3300 -4375 -3266
rect -4341 -3300 -4296 -3266
rect -4434 -3338 -4296 -3300
rect -4434 -3372 -4375 -3338
rect -4341 -3372 -4296 -3338
rect -4434 -3410 -4296 -3372
rect -4434 -3444 -4375 -3410
rect -4341 -3444 -4296 -3410
rect -4434 -3482 -4296 -3444
rect -4434 -3516 -4375 -3482
rect -4341 -3516 -4296 -3482
rect -4434 -3554 -4296 -3516
rect -4434 -3588 -4375 -3554
rect -4341 -3588 -4296 -3554
rect -4434 -3654 -4296 -3588
rect -4125 -2567 -4079 -2533
rect -4045 -2567 -3994 -2533
rect -4125 -2605 -3994 -2567
rect -4125 -2639 -4079 -2605
rect -4045 -2639 -3994 -2605
rect -4125 -2677 -3994 -2639
rect -4125 -2711 -4079 -2677
rect -4045 -2711 -3994 -2677
rect -4125 -2749 -3994 -2711
rect -3792 -2735 -3434 -2402
rect -4125 -2783 -4079 -2749
rect -4045 -2783 -3994 -2749
rect -4125 -2821 -3994 -2783
rect -4125 -2855 -4079 -2821
rect -4045 -2855 -3994 -2821
rect -4125 -2893 -3994 -2855
rect -4125 -2927 -4079 -2893
rect -4045 -2927 -3994 -2893
rect -4125 -2965 -3994 -2927
rect -4125 -2999 -4079 -2965
rect -4045 -2999 -3994 -2965
rect -4125 -3037 -3994 -2999
rect -4125 -3071 -4079 -3037
rect -4045 -3071 -3994 -3037
rect -4125 -3109 -3994 -3071
rect -4125 -3143 -4079 -3109
rect -4045 -3143 -3994 -3109
rect -4125 -3181 -3994 -3143
rect -4125 -3215 -4079 -3181
rect -4045 -3215 -3994 -3181
rect -4125 -3253 -3994 -3215
rect -4125 -3287 -4079 -3253
rect -4045 -3287 -3994 -3253
rect -4125 -3325 -3994 -3287
rect -4125 -3359 -4079 -3325
rect -4045 -3359 -3994 -3325
rect -4125 -3397 -3994 -3359
rect -3792 -3361 -3434 -3028
rect -3253 -3372 -3053 -2255
rect -4125 -3431 -4079 -3397
rect -4045 -3431 -3994 -3397
rect -4125 -3469 -3994 -3431
rect -4125 -3503 -4079 -3469
rect -4045 -3503 -3994 -3469
rect -4125 -3517 -3994 -3503
rect -2853 -3517 -2653 -2426
rect -2453 -3372 -2253 -2255
rect -2053 -3517 -1853 -2426
rect -1653 -3372 -1453 -2255
rect -1253 -3517 -1053 -2426
rect -853 -3372 -653 -2255
rect -453 -3517 -253 -2426
rect -53 -3372 147 -2255
rect 347 -3517 547 -2426
rect 747 -3372 947 -2255
rect 2519 -2364 2589 -437
rect 1147 -3517 1347 -2426
rect 1604 -2434 2589 -2364
rect 2629 -2469 2699 -283
rect 2290 -2503 2402 -2478
rect 2290 -2537 2327 -2503
rect 2361 -2537 2402 -2503
rect 2290 -2575 2402 -2537
rect 2290 -2609 2327 -2575
rect 2361 -2609 2402 -2575
rect 2290 -2647 2402 -2609
rect 2290 -2681 2327 -2647
rect 2361 -2681 2402 -2647
rect 1621 -3043 1979 -2710
rect 2290 -2719 2402 -2681
rect 2290 -2753 2327 -2719
rect 2361 -2753 2402 -2719
rect 2290 -2791 2402 -2753
rect 2290 -2825 2327 -2791
rect 2361 -2825 2402 -2791
rect 2290 -2863 2402 -2825
rect 2290 -2897 2327 -2863
rect 2361 -2897 2402 -2863
rect 2290 -2935 2402 -2897
rect 2290 -2969 2327 -2935
rect 2361 -2969 2402 -2935
rect 2290 -3007 2402 -2969
rect 2290 -3041 2327 -3007
rect 2361 -3041 2402 -3007
rect 2290 -3079 2402 -3041
rect 2290 -3113 2327 -3079
rect 2361 -3113 2402 -3079
rect 2290 -3151 2402 -3113
rect 2290 -3185 2327 -3151
rect 2361 -3185 2402 -3151
rect 2290 -3223 2402 -3185
rect 1598 -3296 2228 -3239
rect 1598 -3412 1631 -3296
rect 2195 -3412 2228 -3296
rect 1598 -3466 2228 -3412
rect 2290 -3257 2327 -3223
rect 2361 -3257 2402 -3223
rect 2290 -3295 2402 -3257
rect 2290 -3329 2327 -3295
rect 2361 -3329 2402 -3295
rect 2290 -3367 2402 -3329
rect 2290 -3401 2327 -3367
rect 2361 -3401 2402 -3367
rect 2290 -3439 2402 -3401
rect 2290 -3473 2327 -3439
rect 2361 -3473 2402 -3439
rect 2290 -3511 2402 -3473
rect 2290 -3517 2327 -3511
rect -4125 -3545 2327 -3517
rect 2361 -3545 2402 -3511
rect -4125 -3548 2402 -3545
rect -4125 -3582 -3970 -3548
rect -3936 -3582 -3898 -3548
rect -3864 -3582 -3826 -3548
rect -3792 -3582 -3754 -3548
rect -3720 -3582 -3682 -3548
rect -3648 -3582 -3610 -3548
rect -3576 -3582 -3538 -3548
rect -3504 -3582 -3466 -3548
rect -3432 -3582 -3394 -3548
rect -3360 -3582 -3322 -3548
rect -3288 -3582 -3250 -3548
rect -3216 -3582 -3178 -3548
rect -3144 -3582 -3106 -3548
rect -3072 -3582 -3034 -3548
rect -3000 -3582 -2962 -3548
rect -2928 -3582 -2890 -3548
rect -2856 -3582 -2818 -3548
rect -2784 -3582 -2746 -3548
rect -2712 -3582 -2674 -3548
rect -2640 -3582 -2602 -3548
rect -2568 -3582 -2530 -3548
rect -2496 -3582 -2458 -3548
rect -2424 -3582 -2386 -3548
rect -2352 -3582 -2314 -3548
rect -2280 -3582 -2242 -3548
rect -2208 -3582 -2170 -3548
rect -2136 -3582 -2098 -3548
rect -2064 -3582 -2026 -3548
rect -1992 -3582 -1954 -3548
rect -1920 -3582 -1882 -3548
rect -1848 -3582 -1810 -3548
rect -1776 -3582 -1738 -3548
rect -1704 -3582 -1666 -3548
rect -1632 -3582 -1594 -3548
rect -1560 -3582 -1522 -3548
rect -1488 -3582 -1450 -3548
rect -1416 -3582 -1378 -3548
rect -1344 -3582 -1306 -3548
rect -1272 -3582 -1234 -3548
rect -1200 -3582 -1162 -3548
rect -1128 -3582 -1090 -3548
rect -1056 -3582 -1018 -3548
rect -984 -3582 -946 -3548
rect -912 -3582 -874 -3548
rect -840 -3582 -802 -3548
rect -768 -3582 -730 -3548
rect -696 -3582 -658 -3548
rect -624 -3582 -586 -3548
rect -552 -3582 -514 -3548
rect -480 -3582 -442 -3548
rect -408 -3582 -370 -3548
rect -336 -3582 -298 -3548
rect -264 -3582 -226 -3548
rect -192 -3582 -154 -3548
rect -120 -3582 -82 -3548
rect -48 -3582 -10 -3548
rect 24 -3582 62 -3548
rect 96 -3582 134 -3548
rect 168 -3582 206 -3548
rect 240 -3582 278 -3548
rect 312 -3582 350 -3548
rect 384 -3582 422 -3548
rect 456 -3582 494 -3548
rect 528 -3582 566 -3548
rect 600 -3582 638 -3548
rect 672 -3582 710 -3548
rect 744 -3582 782 -3548
rect 816 -3582 854 -3548
rect 888 -3582 926 -3548
rect 960 -3582 998 -3548
rect 1032 -3582 1070 -3548
rect 1104 -3582 1142 -3548
rect 1176 -3582 1214 -3548
rect 1248 -3582 1286 -3548
rect 1320 -3582 1358 -3548
rect 1392 -3582 1430 -3548
rect 1464 -3582 1502 -3548
rect 1536 -3582 1574 -3548
rect 1608 -3582 1646 -3548
rect 1680 -3582 1718 -3548
rect 1752 -3582 1790 -3548
rect 1824 -3582 1862 -3548
rect 1896 -3582 1934 -3548
rect 1968 -3582 2006 -3548
rect 2040 -3582 2078 -3548
rect 2112 -3582 2150 -3548
rect 2184 -3582 2222 -3548
rect 2256 -3582 2402 -3548
rect -4125 -3606 2402 -3582
rect 2561 -2500 2699 -2469
rect 2561 -2534 2610 -2500
rect 2644 -2534 2699 -2500
rect 2561 -2572 2699 -2534
rect 2561 -2606 2610 -2572
rect 2644 -2606 2699 -2572
rect 2561 -2644 2699 -2606
rect 2561 -2678 2610 -2644
rect 2644 -2678 2699 -2644
rect 2561 -2716 2699 -2678
rect 2561 -2750 2610 -2716
rect 2644 -2750 2699 -2716
rect 2561 -2788 2699 -2750
rect 2561 -2822 2610 -2788
rect 2644 -2822 2699 -2788
rect 2561 -2860 2699 -2822
rect 2561 -2894 2610 -2860
rect 2644 -2894 2699 -2860
rect 2561 -2932 2699 -2894
rect 2561 -2966 2610 -2932
rect 2644 -2966 2699 -2932
rect 2561 -3004 2699 -2966
rect 2561 -3038 2610 -3004
rect 2644 -3038 2699 -3004
rect 2561 -3076 2699 -3038
rect 2561 -3110 2610 -3076
rect 2644 -3110 2699 -3076
rect 2561 -3148 2699 -3110
rect 2561 -3182 2610 -3148
rect 2644 -3182 2699 -3148
rect 2561 -3231 2699 -3182
rect 2561 -3481 2576 -3231
rect 2682 -3234 2699 -3231
rect 2690 -3286 2699 -3234
rect 2682 -3298 2699 -3286
rect 2690 -3350 2699 -3298
rect 2682 -3362 2699 -3350
rect 2690 -3414 2699 -3362
rect 2682 -3426 2699 -3414
rect 2690 -3478 2699 -3426
rect 2682 -3481 2699 -3478
rect 2561 -3654 2699 -3481
rect -4434 -3696 2699 -3654
rect -4434 -3730 -4371 -3696
rect -4337 -3730 -4299 -3696
rect -4265 -3730 -4227 -3696
rect -4193 -3730 -4155 -3696
rect -4121 -3730 -4083 -3696
rect -4049 -3730 -4011 -3696
rect -3977 -3730 -3939 -3696
rect -3905 -3730 -3867 -3696
rect -3833 -3730 -3795 -3696
rect -3761 -3730 -3723 -3696
rect -3689 -3730 -3651 -3696
rect -3617 -3730 -3579 -3696
rect -3545 -3730 -3507 -3696
rect -3473 -3730 -3435 -3696
rect -3401 -3730 -3363 -3696
rect -3329 -3730 -3291 -3696
rect -3257 -3730 -3219 -3696
rect -3185 -3730 -3147 -3696
rect -3113 -3730 -3075 -3696
rect -3041 -3730 -3003 -3696
rect -2969 -3730 -2931 -3696
rect -2897 -3730 -2859 -3696
rect -2825 -3730 -2787 -3696
rect -2753 -3730 -2715 -3696
rect -2681 -3730 -2643 -3696
rect -2609 -3730 -2571 -3696
rect -2537 -3730 -2499 -3696
rect -2465 -3730 -2427 -3696
rect -2393 -3730 -2355 -3696
rect -2321 -3730 -2283 -3696
rect -2249 -3730 -2211 -3696
rect -2177 -3730 -2139 -3696
rect -2105 -3730 -2067 -3696
rect -2033 -3730 -1995 -3696
rect -1961 -3730 -1923 -3696
rect -1889 -3730 -1851 -3696
rect -1817 -3730 -1779 -3696
rect -1745 -3730 -1707 -3696
rect -1673 -3730 -1635 -3696
rect -1601 -3730 -1563 -3696
rect -1529 -3730 -1491 -3696
rect -1457 -3730 -1419 -3696
rect -1385 -3730 -1347 -3696
rect -1313 -3730 -1275 -3696
rect -1241 -3730 -1203 -3696
rect -1169 -3730 -1131 -3696
rect -1097 -3730 -1059 -3696
rect -1025 -3730 -987 -3696
rect -953 -3730 -915 -3696
rect -881 -3730 -843 -3696
rect -809 -3730 -771 -3696
rect -737 -3730 -699 -3696
rect -665 -3730 -627 -3696
rect -593 -3730 -555 -3696
rect -521 -3730 -483 -3696
rect -449 -3730 -411 -3696
rect -377 -3730 -339 -3696
rect -305 -3730 -267 -3696
rect -233 -3730 -195 -3696
rect -161 -3730 -123 -3696
rect -89 -3730 -51 -3696
rect -17 -3730 21 -3696
rect 55 -3730 93 -3696
rect 127 -3730 165 -3696
rect 199 -3730 237 -3696
rect 271 -3730 309 -3696
rect 343 -3730 381 -3696
rect 415 -3730 453 -3696
rect 487 -3730 525 -3696
rect 559 -3730 597 -3696
rect 631 -3730 669 -3696
rect 703 -3730 741 -3696
rect 775 -3730 813 -3696
rect 847 -3730 885 -3696
rect 919 -3730 957 -3696
rect 991 -3730 1029 -3696
rect 1063 -3730 1101 -3696
rect 1135 -3730 1173 -3696
rect 1207 -3730 1245 -3696
rect 1279 -3730 1317 -3696
rect 1351 -3730 1389 -3696
rect 1423 -3730 1461 -3696
rect 1495 -3730 1533 -3696
rect 1567 -3730 1605 -3696
rect 1639 -3730 1677 -3696
rect 1711 -3730 1749 -3696
rect 1783 -3730 1821 -3696
rect 1855 -3730 1893 -3696
rect 1927 -3730 1965 -3696
rect 1999 -3730 2037 -3696
rect 2071 -3730 2109 -3696
rect 2143 -3730 2181 -3696
rect 2215 -3730 2253 -3696
rect 2287 -3730 2325 -3696
rect 2359 -3730 2397 -3696
rect 2431 -3730 2469 -3696
rect 2503 -3730 2541 -3696
rect 2575 -3730 2613 -3696
rect 2647 -3730 2699 -3696
rect -4434 -3792 2699 -3730
<< via1 >>
rect -4326 6470 2638 6475
rect -4326 6364 -4317 6470
rect -4317 6364 2629 6470
rect 2629 6364 2638 6470
rect -4326 6359 2638 6364
rect -4066 5997 -4014 6049
rect -4002 5997 -3950 6049
rect -3750 5997 -3698 6049
rect -3686 5997 -3634 6049
rect -3434 5997 -3382 6049
rect -3370 5997 -3318 6049
rect -3118 5997 -3066 6049
rect -3054 5997 -3002 6049
rect -2802 5997 -2750 6049
rect -2738 5997 -2686 6049
rect -2486 5997 -2434 6049
rect -2422 5997 -2370 6049
rect -2170 5997 -2118 6049
rect -2106 5997 -2054 6049
rect -1854 5997 -1802 6049
rect -1790 5997 -1738 6049
rect -1538 5997 -1486 6049
rect -1474 5997 -1422 6049
rect -1222 5997 -1170 6049
rect -1158 5997 -1106 6049
rect -906 5997 -854 6049
rect -842 5997 -790 6049
rect -590 5997 -538 6049
rect -526 5997 -474 6049
rect -274 5997 -222 6049
rect -210 5997 -158 6049
rect 42 5997 94 6049
rect 106 5997 158 6049
rect 358 5997 410 6049
rect 422 5997 474 6049
rect 674 5997 726 6049
rect 738 5997 790 6049
rect 990 5997 1042 6049
rect 1054 5997 1106 6049
rect 1306 5997 1358 6049
rect 1370 5997 1422 6049
rect 1622 5997 1674 6049
rect 1686 5997 1738 6049
rect 1938 5997 1990 6049
rect 2002 5997 2054 6049
rect 2254 5997 2306 6049
rect 2318 5997 2370 6049
rect -3908 5872 -3856 5924
rect -3844 5872 -3792 5924
rect -3592 5872 -3540 5924
rect -3528 5872 -3476 5924
rect -3276 5872 -3224 5924
rect -3212 5872 -3160 5924
rect -2960 5872 -2908 5924
rect -2896 5872 -2844 5924
rect -2644 5872 -2592 5924
rect -2580 5872 -2528 5924
rect -2328 5872 -2276 5924
rect -2264 5872 -2212 5924
rect -2012 5872 -1960 5924
rect -1948 5872 -1896 5924
rect -1696 5872 -1644 5924
rect -1632 5872 -1580 5924
rect -1380 5872 -1328 5924
rect -1316 5872 -1264 5924
rect -1064 5872 -1012 5924
rect -1000 5872 -948 5924
rect -748 5872 -696 5924
rect -684 5872 -632 5924
rect -432 5872 -380 5924
rect -368 5872 -316 5924
rect -116 5872 -64 5924
rect -52 5872 0 5924
rect 200 5872 252 5924
rect 264 5872 316 5924
rect 516 5872 568 5924
rect 580 5872 632 5924
rect 832 5872 884 5924
rect 896 5872 948 5924
rect 1148 5872 1200 5924
rect 1212 5872 1264 5924
rect 1464 5872 1516 5924
rect 1528 5872 1580 5924
rect 1780 5872 1832 5924
rect 1844 5872 1896 5924
rect 2096 5872 2148 5924
rect 2160 5872 2212 5924
rect -4066 5557 -4014 5609
rect -4002 5557 -3950 5609
rect -3750 5557 -3698 5609
rect -3686 5557 -3634 5609
rect -3434 5557 -3382 5609
rect -3370 5557 -3318 5609
rect -3118 5557 -3066 5609
rect -3054 5557 -3002 5609
rect -2802 5557 -2750 5609
rect -2738 5557 -2686 5609
rect -2486 5557 -2434 5609
rect -2422 5557 -2370 5609
rect -2170 5557 -2118 5609
rect -2106 5557 -2054 5609
rect -1854 5557 -1802 5609
rect -1790 5557 -1738 5609
rect -1538 5557 -1486 5609
rect -1474 5557 -1422 5609
rect -1222 5557 -1170 5609
rect -1158 5557 -1106 5609
rect -906 5557 -854 5609
rect -842 5557 -790 5609
rect -590 5557 -538 5609
rect -526 5557 -474 5609
rect -274 5557 -222 5609
rect -210 5557 -158 5609
rect 42 5557 94 5609
rect 106 5557 158 5609
rect 358 5557 410 5609
rect 422 5557 474 5609
rect 674 5557 726 5609
rect 738 5557 790 5609
rect 990 5557 1042 5609
rect 1054 5557 1106 5609
rect 1306 5557 1358 5609
rect 1370 5557 1422 5609
rect 1622 5557 1674 5609
rect 1686 5557 1738 5609
rect 1938 5557 1990 5609
rect 2002 5557 2054 5609
rect 2254 5557 2306 5609
rect 2318 5557 2370 5609
rect -3908 5432 -3856 5484
rect -3844 5432 -3792 5484
rect -3592 5432 -3540 5484
rect -3528 5432 -3476 5484
rect -3276 5432 -3224 5484
rect -3212 5432 -3160 5484
rect -2960 5432 -2908 5484
rect -2896 5432 -2844 5484
rect -2644 5432 -2592 5484
rect -2580 5432 -2528 5484
rect -2328 5432 -2276 5484
rect -2264 5432 -2212 5484
rect -2012 5432 -1960 5484
rect -1948 5432 -1896 5484
rect -1696 5432 -1644 5484
rect -1632 5432 -1580 5484
rect -1380 5432 -1328 5484
rect -1316 5432 -1264 5484
rect -1064 5432 -1012 5484
rect -1000 5432 -948 5484
rect -748 5432 -696 5484
rect -684 5432 -632 5484
rect -432 5432 -380 5484
rect -368 5432 -316 5484
rect -116 5432 -64 5484
rect -52 5432 0 5484
rect 200 5432 252 5484
rect 264 5432 316 5484
rect 516 5432 568 5484
rect 580 5432 632 5484
rect 832 5432 884 5484
rect 896 5432 948 5484
rect 1148 5432 1200 5484
rect 1212 5432 1264 5484
rect 1464 5432 1516 5484
rect 1528 5432 1580 5484
rect 1780 5432 1832 5484
rect 1844 5432 1896 5484
rect 2096 5432 2148 5484
rect 2160 5432 2212 5484
rect -4066 5117 -4014 5169
rect -4002 5117 -3950 5169
rect -3750 5117 -3698 5169
rect -3686 5117 -3634 5169
rect -3434 5117 -3382 5169
rect -3370 5117 -3318 5169
rect -3118 5117 -3066 5169
rect -3054 5117 -3002 5169
rect -2802 5117 -2750 5169
rect -2738 5117 -2686 5169
rect -2486 5117 -2434 5169
rect -2422 5117 -2370 5169
rect -2170 5117 -2118 5169
rect -2106 5117 -2054 5169
rect -1854 5117 -1802 5169
rect -1790 5117 -1738 5169
rect -1538 5117 -1486 5169
rect -1474 5117 -1422 5169
rect -1222 5117 -1170 5169
rect -1158 5117 -1106 5169
rect -906 5117 -854 5169
rect -842 5117 -790 5169
rect -590 5117 -538 5169
rect -526 5117 -474 5169
rect -274 5117 -222 5169
rect -210 5117 -158 5169
rect 42 5117 94 5169
rect 106 5117 158 5169
rect 358 5117 410 5169
rect 422 5117 474 5169
rect 674 5117 726 5169
rect 738 5117 790 5169
rect 990 5117 1042 5169
rect 1054 5117 1106 5169
rect 1306 5117 1358 5169
rect 1370 5117 1422 5169
rect 1622 5117 1674 5169
rect 1686 5117 1738 5169
rect 1938 5117 1990 5169
rect 2002 5117 2054 5169
rect 2254 5117 2306 5169
rect 2318 5117 2370 5169
rect -3908 4992 -3856 5044
rect -3844 4992 -3792 5044
rect -3592 4992 -3540 5044
rect -3528 4992 -3476 5044
rect -3276 4992 -3224 5044
rect -3212 4992 -3160 5044
rect -2960 4992 -2908 5044
rect -2896 4992 -2844 5044
rect -2644 4992 -2592 5044
rect -2580 4992 -2528 5044
rect -2328 4992 -2276 5044
rect -2264 4992 -2212 5044
rect -2012 4992 -1960 5044
rect -1948 4992 -1896 5044
rect -1696 4992 -1644 5044
rect -1632 4992 -1580 5044
rect -1380 4992 -1328 5044
rect -1316 4992 -1264 5044
rect -1064 4992 -1012 5044
rect -1000 4992 -948 5044
rect -748 4992 -696 5044
rect -684 4992 -632 5044
rect -432 4992 -380 5044
rect -368 4992 -316 5044
rect -116 4992 -64 5044
rect -52 4992 0 5044
rect 200 4992 252 5044
rect 264 4992 316 5044
rect 516 4992 568 5044
rect 580 4992 632 5044
rect 832 4992 884 5044
rect 896 4992 948 5044
rect 1148 4992 1200 5044
rect 1212 4992 1264 5044
rect 1464 4992 1516 5044
rect 1528 4992 1580 5044
rect 1780 4992 1832 5044
rect 1844 4992 1896 5044
rect 2096 4992 2148 5044
rect 2160 4992 2212 5044
rect -4066 4682 -4014 4734
rect -4002 4682 -3950 4734
rect -3750 4682 -3698 4734
rect -3686 4682 -3634 4734
rect -3434 4682 -3382 4734
rect -3370 4682 -3318 4734
rect -3118 4682 -3066 4734
rect -3054 4682 -3002 4734
rect -2802 4682 -2750 4734
rect -2738 4682 -2686 4734
rect -2486 4682 -2434 4734
rect -2422 4682 -2370 4734
rect -2170 4682 -2118 4734
rect -2106 4682 -2054 4734
rect -1854 4682 -1802 4734
rect -1790 4682 -1738 4734
rect -1538 4682 -1486 4734
rect -1474 4682 -1422 4734
rect -1222 4682 -1170 4734
rect -1158 4682 -1106 4734
rect -906 4682 -854 4734
rect -842 4682 -790 4734
rect -590 4682 -538 4734
rect -526 4682 -474 4734
rect -274 4682 -222 4734
rect -210 4682 -158 4734
rect 42 4682 94 4734
rect 106 4682 158 4734
rect 358 4682 410 4734
rect 422 4682 474 4734
rect 674 4682 726 4734
rect 738 4682 790 4734
rect 990 4682 1042 4734
rect 1054 4682 1106 4734
rect 1306 4682 1358 4734
rect 1370 4682 1422 4734
rect 1622 4682 1674 4734
rect 1686 4682 1738 4734
rect 1938 4682 1990 4734
rect 2002 4682 2054 4734
rect 2254 4682 2306 4734
rect 2318 4682 2370 4734
rect -3908 4557 -3856 4609
rect -3844 4557 -3792 4609
rect -3592 4557 -3540 4609
rect -3528 4557 -3476 4609
rect -3276 4557 -3224 4609
rect -3212 4557 -3160 4609
rect -2960 4557 -2908 4609
rect -2896 4557 -2844 4609
rect -2644 4557 -2592 4609
rect -2580 4557 -2528 4609
rect -2328 4557 -2276 4609
rect -2264 4557 -2212 4609
rect -2012 4557 -1960 4609
rect -1948 4557 -1896 4609
rect -1696 4557 -1644 4609
rect -1632 4557 -1580 4609
rect -1380 4557 -1328 4609
rect -1316 4557 -1264 4609
rect -1064 4557 -1012 4609
rect -1000 4557 -948 4609
rect -748 4557 -696 4609
rect -684 4557 -632 4609
rect -432 4557 -380 4609
rect -368 4557 -316 4609
rect -116 4557 -64 4609
rect -52 4557 0 4609
rect 200 4557 252 4609
rect 264 4557 316 4609
rect 516 4557 568 4609
rect 580 4557 632 4609
rect 832 4557 884 4609
rect 896 4557 948 4609
rect 1148 4557 1200 4609
rect 1212 4557 1264 4609
rect 1464 4557 1516 4609
rect 1528 4557 1580 4609
rect 1780 4557 1832 4609
rect 1844 4557 1896 4609
rect 2096 4557 2148 4609
rect 2160 4557 2212 4609
rect -4066 4257 -4014 4309
rect -4002 4257 -3950 4309
rect -3750 4257 -3698 4309
rect -3686 4257 -3634 4309
rect -3434 4257 -3382 4309
rect -3370 4257 -3318 4309
rect -3118 4257 -3066 4309
rect -3054 4257 -3002 4309
rect -2802 4257 -2750 4309
rect -2738 4257 -2686 4309
rect -2486 4257 -2434 4309
rect -2422 4257 -2370 4309
rect -2170 4257 -2118 4309
rect -2106 4257 -2054 4309
rect -1854 4257 -1802 4309
rect -1790 4257 -1738 4309
rect -1538 4257 -1486 4309
rect -1474 4257 -1422 4309
rect -1222 4257 -1170 4309
rect -1158 4257 -1106 4309
rect -906 4257 -854 4309
rect -842 4257 -790 4309
rect -590 4257 -538 4309
rect -526 4257 -474 4309
rect -274 4257 -222 4309
rect -210 4257 -158 4309
rect 42 4257 94 4309
rect 106 4257 158 4309
rect 358 4257 410 4309
rect 422 4257 474 4309
rect 674 4257 726 4309
rect 738 4257 790 4309
rect 990 4257 1042 4309
rect 1054 4257 1106 4309
rect 1306 4257 1358 4309
rect 1370 4257 1422 4309
rect 1622 4257 1674 4309
rect 1686 4257 1738 4309
rect 1938 4257 1990 4309
rect 2002 4257 2054 4309
rect 2254 4257 2306 4309
rect 2318 4257 2370 4309
rect -3908 4132 -3856 4184
rect -3844 4132 -3792 4184
rect -3592 4132 -3540 4184
rect -3528 4132 -3476 4184
rect -3276 4132 -3224 4184
rect -3212 4132 -3160 4184
rect -2960 4132 -2908 4184
rect -2896 4132 -2844 4184
rect -2644 4132 -2592 4184
rect -2580 4132 -2528 4184
rect -2328 4132 -2276 4184
rect -2264 4132 -2212 4184
rect -2012 4132 -1960 4184
rect -1948 4132 -1896 4184
rect -1696 4132 -1644 4184
rect -1632 4132 -1580 4184
rect -1380 4132 -1328 4184
rect -1316 4132 -1264 4184
rect -1064 4132 -1012 4184
rect -1000 4132 -948 4184
rect -748 4132 -696 4184
rect -684 4132 -632 4184
rect -432 4132 -380 4184
rect -368 4132 -316 4184
rect -116 4132 -64 4184
rect -52 4132 0 4184
rect 200 4132 252 4184
rect 264 4132 316 4184
rect 516 4132 568 4184
rect 580 4132 632 4184
rect 832 4132 884 4184
rect 896 4132 948 4184
rect 1148 4132 1200 4184
rect 1212 4132 1264 4184
rect 1464 4132 1516 4184
rect 1528 4132 1580 4184
rect 1780 4132 1832 4184
rect 1844 4132 1896 4184
rect 2096 4132 2148 4184
rect 2160 4132 2212 4184
rect -4110 3926 -4058 3937
rect -4046 3926 -3994 3937
rect -3982 3926 -3930 3937
rect -3918 3926 -3866 3937
rect -3854 3926 -3802 3937
rect -4110 3892 -4076 3926
rect -4076 3892 -4058 3926
rect -4046 3892 -4042 3926
rect -4042 3892 -4004 3926
rect -4004 3892 -3994 3926
rect -3982 3892 -3970 3926
rect -3970 3892 -3932 3926
rect -3932 3892 -3930 3926
rect -3918 3892 -3898 3926
rect -3898 3892 -3866 3926
rect -3854 3892 -3826 3926
rect -3826 3892 -3802 3926
rect -4110 3885 -4058 3892
rect -4046 3885 -3994 3892
rect -3982 3885 -3930 3892
rect -3918 3885 -3866 3892
rect -3854 3885 -3802 3892
rect -3790 3926 -3738 3937
rect -3790 3892 -3788 3926
rect -3788 3892 -3754 3926
rect -3754 3892 -3738 3926
rect -3790 3885 -3738 3892
rect -3726 3926 -3674 3937
rect -3726 3892 -3716 3926
rect -3716 3892 -3682 3926
rect -3682 3892 -3674 3926
rect -3726 3885 -3674 3892
rect -3662 3926 -3610 3937
rect -3662 3892 -3644 3926
rect -3644 3892 -3610 3926
rect -3662 3885 -3610 3892
rect -3598 3926 -3546 3937
rect -3534 3926 -3482 3937
rect -3470 3926 -3418 3937
rect -3406 3926 -3354 3937
rect -3342 3926 -3290 3937
rect -3278 3926 -3226 3937
rect -3598 3892 -3572 3926
rect -3572 3892 -3546 3926
rect -3534 3892 -3500 3926
rect -3500 3892 -3482 3926
rect -3470 3892 -3466 3926
rect -3466 3892 -3428 3926
rect -3428 3892 -3418 3926
rect -3406 3892 -3394 3926
rect -3394 3892 -3356 3926
rect -3356 3892 -3354 3926
rect -3342 3892 -3322 3926
rect -3322 3892 -3290 3926
rect -3278 3892 -3250 3926
rect -3250 3892 -3226 3926
rect -3598 3885 -3546 3892
rect -3534 3885 -3482 3892
rect -3470 3885 -3418 3892
rect -3406 3885 -3354 3892
rect -3342 3885 -3290 3892
rect -3278 3885 -3226 3892
rect -3214 3926 -3162 3937
rect -3214 3892 -3212 3926
rect -3212 3892 -3178 3926
rect -3178 3892 -3162 3926
rect -3214 3885 -3162 3892
rect -3150 3926 -3098 3937
rect -3150 3892 -3140 3926
rect -3140 3892 -3106 3926
rect -3106 3892 -3098 3926
rect -3150 3885 -3098 3892
rect -3086 3926 -3034 3937
rect -3086 3892 -3068 3926
rect -3068 3892 -3034 3926
rect -3086 3885 -3034 3892
rect -3022 3926 -2970 3937
rect -2958 3926 -2906 3937
rect -2894 3926 -2842 3937
rect -2830 3926 -2778 3937
rect -2766 3926 -2714 3937
rect -2702 3926 -2650 3937
rect -3022 3892 -2996 3926
rect -2996 3892 -2970 3926
rect -2958 3892 -2924 3926
rect -2924 3892 -2906 3926
rect -2894 3892 -2890 3926
rect -2890 3892 -2852 3926
rect -2852 3892 -2842 3926
rect -2830 3892 -2818 3926
rect -2818 3892 -2780 3926
rect -2780 3892 -2778 3926
rect -2766 3892 -2746 3926
rect -2746 3892 -2714 3926
rect -2702 3892 -2674 3926
rect -2674 3892 -2650 3926
rect -3022 3885 -2970 3892
rect -2958 3885 -2906 3892
rect -2894 3885 -2842 3892
rect -2830 3885 -2778 3892
rect -2766 3885 -2714 3892
rect -2702 3885 -2650 3892
rect -2638 3926 -2586 3937
rect -2638 3892 -2636 3926
rect -2636 3892 -2602 3926
rect -2602 3892 -2586 3926
rect -2638 3885 -2586 3892
rect -2574 3926 -2522 3937
rect -2574 3892 -2564 3926
rect -2564 3892 -2530 3926
rect -2530 3892 -2522 3926
rect -2574 3885 -2522 3892
rect -2510 3926 -2458 3937
rect -2510 3892 -2492 3926
rect -2492 3892 -2458 3926
rect -2510 3885 -2458 3892
rect -2446 3926 -2394 3937
rect -2382 3926 -2330 3937
rect -2318 3926 -2266 3937
rect -2254 3926 -2202 3937
rect -2190 3926 -2138 3937
rect -2126 3926 -2074 3937
rect -2446 3892 -2420 3926
rect -2420 3892 -2394 3926
rect -2382 3892 -2348 3926
rect -2348 3892 -2330 3926
rect -2318 3892 -2314 3926
rect -2314 3892 -2276 3926
rect -2276 3892 -2266 3926
rect -2254 3892 -2242 3926
rect -2242 3892 -2204 3926
rect -2204 3892 -2202 3926
rect -2190 3892 -2170 3926
rect -2170 3892 -2138 3926
rect -2126 3892 -2098 3926
rect -2098 3892 -2074 3926
rect -2446 3885 -2394 3892
rect -2382 3885 -2330 3892
rect -2318 3885 -2266 3892
rect -2254 3885 -2202 3892
rect -2190 3885 -2138 3892
rect -2126 3885 -2074 3892
rect -2062 3926 -2010 3937
rect -2062 3892 -2060 3926
rect -2060 3892 -2026 3926
rect -2026 3892 -2010 3926
rect -2062 3885 -2010 3892
rect -1998 3926 -1946 3937
rect -1998 3892 -1988 3926
rect -1988 3892 -1954 3926
rect -1954 3892 -1946 3926
rect -1998 3885 -1946 3892
rect -1934 3926 -1882 3937
rect -1934 3892 -1916 3926
rect -1916 3892 -1882 3926
rect -1934 3885 -1882 3892
rect -1870 3926 -1818 3937
rect -1806 3926 -1754 3937
rect -1742 3926 -1690 3937
rect -1678 3926 -1626 3937
rect -1614 3926 -1562 3937
rect -1550 3926 -1498 3937
rect -1870 3892 -1844 3926
rect -1844 3892 -1818 3926
rect -1806 3892 -1772 3926
rect -1772 3892 -1754 3926
rect -1742 3892 -1738 3926
rect -1738 3892 -1700 3926
rect -1700 3892 -1690 3926
rect -1678 3892 -1666 3926
rect -1666 3892 -1628 3926
rect -1628 3892 -1626 3926
rect -1614 3892 -1594 3926
rect -1594 3892 -1562 3926
rect -1550 3892 -1522 3926
rect -1522 3892 -1498 3926
rect -1870 3885 -1818 3892
rect -1806 3885 -1754 3892
rect -1742 3885 -1690 3892
rect -1678 3885 -1626 3892
rect -1614 3885 -1562 3892
rect -1550 3885 -1498 3892
rect -1486 3926 -1434 3937
rect -1486 3892 -1484 3926
rect -1484 3892 -1450 3926
rect -1450 3892 -1434 3926
rect -1486 3885 -1434 3892
rect -1422 3926 -1370 3937
rect -1422 3892 -1412 3926
rect -1412 3892 -1378 3926
rect -1378 3892 -1370 3926
rect -1422 3885 -1370 3892
rect -1358 3926 -1306 3937
rect -1358 3892 -1340 3926
rect -1340 3892 -1306 3926
rect -1358 3885 -1306 3892
rect -1294 3926 -1242 3937
rect -1230 3926 -1178 3937
rect -1166 3926 -1114 3937
rect -1102 3926 -1050 3937
rect -1038 3926 -986 3937
rect -974 3926 -922 3937
rect -1294 3892 -1268 3926
rect -1268 3892 -1242 3926
rect -1230 3892 -1196 3926
rect -1196 3892 -1178 3926
rect -1166 3892 -1162 3926
rect -1162 3892 -1124 3926
rect -1124 3892 -1114 3926
rect -1102 3892 -1090 3926
rect -1090 3892 -1052 3926
rect -1052 3892 -1050 3926
rect -1038 3892 -1018 3926
rect -1018 3892 -986 3926
rect -974 3892 -946 3926
rect -946 3892 -922 3926
rect -1294 3885 -1242 3892
rect -1230 3885 -1178 3892
rect -1166 3885 -1114 3892
rect -1102 3885 -1050 3892
rect -1038 3885 -986 3892
rect -974 3885 -922 3892
rect -910 3926 -858 3937
rect -910 3892 -908 3926
rect -908 3892 -874 3926
rect -874 3892 -858 3926
rect -910 3885 -858 3892
rect -846 3926 -794 3937
rect -846 3892 -836 3926
rect -836 3892 -802 3926
rect -802 3892 -794 3926
rect -846 3885 -794 3892
rect -782 3926 -730 3937
rect -782 3892 -764 3926
rect -764 3892 -730 3926
rect -782 3885 -730 3892
rect -718 3926 -666 3937
rect -654 3926 -602 3937
rect -590 3926 -538 3937
rect -526 3926 -474 3937
rect -462 3926 -410 3937
rect -398 3926 -346 3937
rect -718 3892 -692 3926
rect -692 3892 -666 3926
rect -654 3892 -620 3926
rect -620 3892 -602 3926
rect -590 3892 -586 3926
rect -586 3892 -548 3926
rect -548 3892 -538 3926
rect -526 3892 -514 3926
rect -514 3892 -476 3926
rect -476 3892 -474 3926
rect -462 3892 -442 3926
rect -442 3892 -410 3926
rect -398 3892 -370 3926
rect -370 3892 -346 3926
rect -718 3885 -666 3892
rect -654 3885 -602 3892
rect -590 3885 -538 3892
rect -526 3885 -474 3892
rect -462 3885 -410 3892
rect -398 3885 -346 3892
rect -334 3926 -282 3937
rect -334 3892 -332 3926
rect -332 3892 -298 3926
rect -298 3892 -282 3926
rect -334 3885 -282 3892
rect -270 3926 -218 3937
rect -270 3892 -260 3926
rect -260 3892 -226 3926
rect -226 3892 -218 3926
rect -270 3885 -218 3892
rect -206 3926 -154 3937
rect -206 3892 -188 3926
rect -188 3892 -154 3926
rect -206 3885 -154 3892
rect -142 3926 -90 3937
rect -78 3926 -26 3937
rect -14 3926 38 3937
rect 50 3926 102 3937
rect 114 3926 166 3937
rect 178 3926 230 3937
rect -142 3892 -116 3926
rect -116 3892 -90 3926
rect -78 3892 -44 3926
rect -44 3892 -26 3926
rect -14 3892 -10 3926
rect -10 3892 28 3926
rect 28 3892 38 3926
rect 50 3892 62 3926
rect 62 3892 100 3926
rect 100 3892 102 3926
rect 114 3892 134 3926
rect 134 3892 166 3926
rect 178 3892 206 3926
rect 206 3892 230 3926
rect -142 3885 -90 3892
rect -78 3885 -26 3892
rect -14 3885 38 3892
rect 50 3885 102 3892
rect 114 3885 166 3892
rect 178 3885 230 3892
rect 242 3926 294 3937
rect 242 3892 244 3926
rect 244 3892 278 3926
rect 278 3892 294 3926
rect 242 3885 294 3892
rect 306 3926 358 3937
rect 306 3892 316 3926
rect 316 3892 350 3926
rect 350 3892 358 3926
rect 306 3885 358 3892
rect 370 3926 422 3937
rect 370 3892 388 3926
rect 388 3892 422 3926
rect 370 3885 422 3892
rect 434 3926 486 3937
rect 498 3926 550 3937
rect 562 3926 614 3937
rect 626 3926 678 3937
rect 690 3926 742 3937
rect 754 3926 806 3937
rect 434 3892 460 3926
rect 460 3892 486 3926
rect 498 3892 532 3926
rect 532 3892 550 3926
rect 562 3892 566 3926
rect 566 3892 604 3926
rect 604 3892 614 3926
rect 626 3892 638 3926
rect 638 3892 676 3926
rect 676 3892 678 3926
rect 690 3892 710 3926
rect 710 3892 742 3926
rect 754 3892 782 3926
rect 782 3892 806 3926
rect 434 3885 486 3892
rect 498 3885 550 3892
rect 562 3885 614 3892
rect 626 3885 678 3892
rect 690 3885 742 3892
rect 754 3885 806 3892
rect 818 3926 870 3937
rect 818 3892 820 3926
rect 820 3892 854 3926
rect 854 3892 870 3926
rect 818 3885 870 3892
rect 882 3926 934 3937
rect 882 3892 892 3926
rect 892 3892 926 3926
rect 926 3892 934 3926
rect 882 3885 934 3892
rect 946 3926 998 3937
rect 946 3892 964 3926
rect 964 3892 998 3926
rect 946 3885 998 3892
rect 1010 3926 1062 3937
rect 1074 3926 1126 3937
rect 1138 3926 1190 3937
rect 1202 3926 1254 3937
rect 1266 3926 1318 3937
rect 1330 3926 1382 3937
rect 1010 3892 1036 3926
rect 1036 3892 1062 3926
rect 1074 3892 1108 3926
rect 1108 3892 1126 3926
rect 1138 3892 1142 3926
rect 1142 3892 1180 3926
rect 1180 3892 1190 3926
rect 1202 3892 1214 3926
rect 1214 3892 1252 3926
rect 1252 3892 1254 3926
rect 1266 3892 1286 3926
rect 1286 3892 1318 3926
rect 1330 3892 1358 3926
rect 1358 3892 1382 3926
rect 1010 3885 1062 3892
rect 1074 3885 1126 3892
rect 1138 3885 1190 3892
rect 1202 3885 1254 3892
rect 1266 3885 1318 3892
rect 1330 3885 1382 3892
rect 1394 3926 1446 3937
rect 1394 3892 1396 3926
rect 1396 3892 1430 3926
rect 1430 3892 1446 3926
rect 1394 3885 1446 3892
rect 1458 3926 1510 3937
rect 1458 3892 1468 3926
rect 1468 3892 1502 3926
rect 1502 3892 1510 3926
rect 1458 3885 1510 3892
rect 1522 3926 1574 3937
rect 1522 3892 1540 3926
rect 1540 3892 1574 3926
rect 1522 3885 1574 3892
rect 1586 3926 1638 3937
rect 1650 3926 1702 3937
rect 1714 3926 1766 3937
rect 1778 3926 1830 3937
rect 1842 3926 1894 3937
rect 1906 3926 1958 3937
rect 1586 3892 1612 3926
rect 1612 3892 1638 3926
rect 1650 3892 1684 3926
rect 1684 3892 1702 3926
rect 1714 3892 1718 3926
rect 1718 3892 1756 3926
rect 1756 3892 1766 3926
rect 1778 3892 1790 3926
rect 1790 3892 1828 3926
rect 1828 3892 1830 3926
rect 1842 3892 1862 3926
rect 1862 3892 1894 3926
rect 1906 3892 1934 3926
rect 1934 3892 1958 3926
rect 1586 3885 1638 3892
rect 1650 3885 1702 3892
rect 1714 3885 1766 3892
rect 1778 3885 1830 3892
rect 1842 3885 1894 3892
rect 1906 3885 1958 3892
rect 1970 3926 2022 3937
rect 1970 3892 1972 3926
rect 1972 3892 2006 3926
rect 2006 3892 2022 3926
rect 1970 3885 2022 3892
rect 2034 3926 2086 3937
rect 2034 3892 2044 3926
rect 2044 3892 2078 3926
rect 2078 3892 2086 3926
rect 2034 3885 2086 3892
rect 2098 3926 2150 3937
rect 2098 3892 2116 3926
rect 2116 3892 2150 3926
rect 2098 3885 2150 3892
rect 2162 3926 2214 3937
rect 2226 3926 2278 3937
rect 2290 3926 2342 3937
rect 2162 3892 2188 3926
rect 2188 3892 2214 3926
rect 2226 3892 2260 3926
rect 2260 3892 2278 3926
rect 2290 3892 2294 3926
rect 2294 3892 2332 3926
rect 2332 3892 2342 3926
rect 2162 3885 2214 3892
rect 2226 3885 2278 3892
rect 2290 3885 2342 3892
rect -4066 3637 -4014 3689
rect -4002 3637 -3950 3689
rect -3750 3637 -3698 3689
rect -3686 3637 -3634 3689
rect -3434 3637 -3382 3689
rect -3370 3637 -3318 3689
rect -3118 3637 -3066 3689
rect -3054 3637 -3002 3689
rect -2802 3637 -2750 3689
rect -2738 3637 -2686 3689
rect -2486 3637 -2434 3689
rect -2422 3637 -2370 3689
rect -2170 3637 -2118 3689
rect -2106 3637 -2054 3689
rect -1854 3637 -1802 3689
rect -1790 3637 -1738 3689
rect -1538 3637 -1486 3689
rect -1474 3637 -1422 3689
rect -1222 3637 -1170 3689
rect -1158 3637 -1106 3689
rect -906 3637 -854 3689
rect -842 3637 -790 3689
rect -590 3637 -538 3689
rect -526 3637 -474 3689
rect -274 3637 -222 3689
rect -210 3637 -158 3689
rect 42 3637 94 3689
rect 106 3637 158 3689
rect 358 3637 410 3689
rect 422 3637 474 3689
rect 674 3637 726 3689
rect 738 3637 790 3689
rect 990 3637 1042 3689
rect 1054 3637 1106 3689
rect 1306 3637 1358 3689
rect 1370 3637 1422 3689
rect 1622 3637 1674 3689
rect 1686 3637 1738 3689
rect 1938 3637 1990 3689
rect 2002 3637 2054 3689
rect 2254 3637 2306 3689
rect 2318 3637 2370 3689
rect -3908 3512 -3856 3564
rect -3844 3512 -3792 3564
rect -3592 3512 -3540 3564
rect -3528 3512 -3476 3564
rect -3276 3512 -3224 3564
rect -3212 3512 -3160 3564
rect -2960 3512 -2908 3564
rect -2896 3512 -2844 3564
rect -2644 3512 -2592 3564
rect -2580 3512 -2528 3564
rect -2328 3512 -2276 3564
rect -2264 3512 -2212 3564
rect -2012 3512 -1960 3564
rect -1948 3512 -1896 3564
rect -1696 3512 -1644 3564
rect -1632 3512 -1580 3564
rect -1380 3512 -1328 3564
rect -1316 3512 -1264 3564
rect -1064 3512 -1012 3564
rect -1000 3512 -948 3564
rect -748 3512 -696 3564
rect -684 3512 -632 3564
rect -432 3512 -380 3564
rect -368 3512 -316 3564
rect -116 3512 -64 3564
rect -52 3512 0 3564
rect 200 3512 252 3564
rect 264 3512 316 3564
rect 516 3512 568 3564
rect 580 3512 632 3564
rect 832 3512 884 3564
rect 896 3512 948 3564
rect 1148 3512 1200 3564
rect 1212 3512 1264 3564
rect 1464 3512 1516 3564
rect 1528 3512 1580 3564
rect 1780 3512 1832 3564
rect 1844 3512 1896 3564
rect 2096 3512 2148 3564
rect 2160 3512 2212 3564
rect -4066 3202 -4014 3254
rect -4002 3202 -3950 3254
rect -3750 3202 -3698 3254
rect -3686 3202 -3634 3254
rect -3434 3202 -3382 3254
rect -3370 3202 -3318 3254
rect -3118 3202 -3066 3254
rect -3054 3202 -3002 3254
rect -2802 3202 -2750 3254
rect -2738 3202 -2686 3254
rect -2486 3202 -2434 3254
rect -2422 3202 -2370 3254
rect -2170 3202 -2118 3254
rect -2106 3202 -2054 3254
rect -1854 3202 -1802 3254
rect -1790 3202 -1738 3254
rect -1538 3202 -1486 3254
rect -1474 3202 -1422 3254
rect -1222 3202 -1170 3254
rect -1158 3202 -1106 3254
rect -906 3202 -854 3254
rect -842 3202 -790 3254
rect -590 3202 -538 3254
rect -526 3202 -474 3254
rect -274 3202 -222 3254
rect -210 3202 -158 3254
rect 42 3202 94 3254
rect 106 3202 158 3254
rect 358 3202 410 3254
rect 422 3202 474 3254
rect 674 3202 726 3254
rect 738 3202 790 3254
rect 990 3202 1042 3254
rect 1054 3202 1106 3254
rect 1306 3202 1358 3254
rect 1370 3202 1422 3254
rect 1622 3202 1674 3254
rect 1686 3202 1738 3254
rect 1938 3202 1990 3254
rect 2002 3202 2054 3254
rect 2254 3202 2306 3254
rect 2318 3202 2370 3254
rect -3908 3077 -3856 3129
rect -3844 3077 -3792 3129
rect -3592 3077 -3540 3129
rect -3528 3077 -3476 3129
rect -3276 3077 -3224 3129
rect -3212 3077 -3160 3129
rect -2960 3077 -2908 3129
rect -2896 3077 -2844 3129
rect -2644 3077 -2592 3129
rect -2580 3077 -2528 3129
rect -2328 3077 -2276 3129
rect -2264 3077 -2212 3129
rect -2012 3077 -1960 3129
rect -1948 3077 -1896 3129
rect -1696 3077 -1644 3129
rect -1632 3077 -1580 3129
rect -1380 3077 -1328 3129
rect -1316 3077 -1264 3129
rect -1064 3077 -1012 3129
rect -1000 3077 -948 3129
rect -748 3077 -696 3129
rect -684 3077 -632 3129
rect -432 3077 -380 3129
rect -368 3077 -316 3129
rect -116 3077 -64 3129
rect -52 3077 0 3129
rect 200 3077 252 3129
rect 264 3077 316 3129
rect 516 3077 568 3129
rect 580 3077 632 3129
rect 832 3077 884 3129
rect 896 3077 948 3129
rect 1148 3077 1200 3129
rect 1212 3077 1264 3129
rect 1464 3077 1516 3129
rect 1528 3077 1580 3129
rect 1780 3077 1832 3129
rect 1844 3077 1896 3129
rect 2096 3077 2148 3129
rect 2160 3077 2212 3129
rect -4066 2767 -4014 2819
rect -4002 2767 -3950 2819
rect -3750 2767 -3698 2819
rect -3686 2767 -3634 2819
rect -3434 2767 -3382 2819
rect -3370 2767 -3318 2819
rect -3118 2767 -3066 2819
rect -3054 2767 -3002 2819
rect -2802 2767 -2750 2819
rect -2738 2767 -2686 2819
rect -2486 2767 -2434 2819
rect -2422 2767 -2370 2819
rect -2170 2767 -2118 2819
rect -2106 2767 -2054 2819
rect -1854 2767 -1802 2819
rect -1790 2767 -1738 2819
rect -1538 2767 -1486 2819
rect -1474 2767 -1422 2819
rect -1222 2767 -1170 2819
rect -1158 2767 -1106 2819
rect -906 2767 -854 2819
rect -842 2767 -790 2819
rect -590 2767 -538 2819
rect -526 2767 -474 2819
rect -274 2767 -222 2819
rect -210 2767 -158 2819
rect 42 2767 94 2819
rect 106 2767 158 2819
rect 358 2767 410 2819
rect 422 2767 474 2819
rect 674 2767 726 2819
rect 738 2767 790 2819
rect 990 2767 1042 2819
rect 1054 2767 1106 2819
rect 1306 2767 1358 2819
rect 1370 2767 1422 2819
rect 1622 2767 1674 2819
rect 1686 2767 1738 2819
rect 1938 2767 1990 2819
rect 2002 2767 2054 2819
rect 2254 2767 2306 2819
rect 2318 2767 2370 2819
rect -3908 2642 -3856 2694
rect -3844 2642 -3792 2694
rect -3592 2642 -3540 2694
rect -3528 2642 -3476 2694
rect -3276 2642 -3224 2694
rect -3212 2642 -3160 2694
rect -2960 2642 -2908 2694
rect -2896 2642 -2844 2694
rect -2644 2642 -2592 2694
rect -2580 2642 -2528 2694
rect -2328 2642 -2276 2694
rect -2264 2642 -2212 2694
rect -2012 2642 -1960 2694
rect -1948 2642 -1896 2694
rect -1696 2642 -1644 2694
rect -1632 2642 -1580 2694
rect -1380 2642 -1328 2694
rect -1316 2642 -1264 2694
rect -1064 2642 -1012 2694
rect -1000 2642 -948 2694
rect -748 2642 -696 2694
rect -684 2642 -632 2694
rect -432 2642 -380 2694
rect -368 2642 -316 2694
rect -116 2642 -64 2694
rect -52 2642 0 2694
rect 200 2642 252 2694
rect 264 2642 316 2694
rect 516 2642 568 2694
rect 580 2642 632 2694
rect 832 2642 884 2694
rect 896 2642 948 2694
rect 1148 2642 1200 2694
rect 1212 2642 1264 2694
rect 1464 2642 1516 2694
rect 1528 2642 1580 2694
rect 1780 2642 1832 2694
rect 1844 2642 1896 2694
rect 2096 2642 2148 2694
rect 2160 2642 2212 2694
rect -4066 2332 -4014 2384
rect -4002 2332 -3950 2384
rect -3750 2332 -3698 2384
rect -3686 2332 -3634 2384
rect -3434 2332 -3382 2384
rect -3370 2332 -3318 2384
rect -3118 2332 -3066 2384
rect -3054 2332 -3002 2384
rect -2802 2332 -2750 2384
rect -2738 2332 -2686 2384
rect -2486 2332 -2434 2384
rect -2422 2332 -2370 2384
rect -2170 2332 -2118 2384
rect -2106 2332 -2054 2384
rect -1854 2332 -1802 2384
rect -1790 2332 -1738 2384
rect -1538 2332 -1486 2384
rect -1474 2332 -1422 2384
rect -1222 2332 -1170 2384
rect -1158 2332 -1106 2384
rect -906 2332 -854 2384
rect -842 2332 -790 2384
rect -590 2332 -538 2384
rect -526 2332 -474 2384
rect -274 2332 -222 2384
rect -210 2332 -158 2384
rect 42 2332 94 2384
rect 106 2332 158 2384
rect 358 2332 410 2384
rect 422 2332 474 2384
rect 674 2332 726 2384
rect 738 2332 790 2384
rect 990 2332 1042 2384
rect 1054 2332 1106 2384
rect 1306 2332 1358 2384
rect 1370 2332 1422 2384
rect 1622 2332 1674 2384
rect 1686 2332 1738 2384
rect 1938 2332 1990 2384
rect 2002 2332 2054 2384
rect 2254 2332 2306 2384
rect 2318 2332 2370 2384
rect -3908 2207 -3856 2259
rect -3844 2207 -3792 2259
rect -3592 2207 -3540 2259
rect -3528 2207 -3476 2259
rect -3276 2207 -3224 2259
rect -3212 2207 -3160 2259
rect -2960 2207 -2908 2259
rect -2896 2207 -2844 2259
rect -2644 2207 -2592 2259
rect -2580 2207 -2528 2259
rect -2328 2207 -2276 2259
rect -2264 2207 -2212 2259
rect -2012 2207 -1960 2259
rect -1948 2207 -1896 2259
rect -1696 2207 -1644 2259
rect -1632 2207 -1580 2259
rect -1380 2207 -1328 2259
rect -1316 2207 -1264 2259
rect -1064 2207 -1012 2259
rect -1000 2207 -948 2259
rect -748 2207 -696 2259
rect -684 2207 -632 2259
rect -432 2207 -380 2259
rect -368 2207 -316 2259
rect -116 2207 -64 2259
rect -52 2207 0 2259
rect 200 2207 252 2259
rect 264 2207 316 2259
rect 516 2207 568 2259
rect 580 2207 632 2259
rect 832 2207 884 2259
rect 896 2207 948 2259
rect 1148 2207 1200 2259
rect 1212 2207 1264 2259
rect 1464 2207 1516 2259
rect 1528 2207 1580 2259
rect 1780 2207 1832 2259
rect 1844 2207 1896 2259
rect 2096 2207 2148 2259
rect 2160 2207 2212 2259
rect -4066 1897 -4014 1949
rect -4002 1897 -3950 1949
rect -3750 1897 -3698 1949
rect -3686 1897 -3634 1949
rect -3434 1897 -3382 1949
rect -3370 1897 -3318 1949
rect -3118 1897 -3066 1949
rect -3054 1897 -3002 1949
rect -2802 1897 -2750 1949
rect -2738 1897 -2686 1949
rect -2486 1897 -2434 1949
rect -2422 1897 -2370 1949
rect -2170 1897 -2118 1949
rect -2106 1897 -2054 1949
rect -1854 1897 -1802 1949
rect -1790 1897 -1738 1949
rect -1538 1897 -1486 1949
rect -1474 1897 -1422 1949
rect -1222 1897 -1170 1949
rect -1158 1897 -1106 1949
rect -906 1897 -854 1949
rect -842 1897 -790 1949
rect -590 1897 -538 1949
rect -526 1897 -474 1949
rect -274 1897 -222 1949
rect -210 1897 -158 1949
rect 42 1897 94 1949
rect 106 1897 158 1949
rect 358 1897 410 1949
rect 422 1897 474 1949
rect 674 1897 726 1949
rect 738 1897 790 1949
rect 990 1897 1042 1949
rect 1054 1897 1106 1949
rect 1306 1897 1358 1949
rect 1370 1897 1422 1949
rect 1622 1897 1674 1949
rect 1686 1897 1738 1949
rect 1938 1897 1990 1949
rect 2002 1897 2054 1949
rect 2254 1897 2306 1949
rect 2318 1897 2370 1949
rect -3908 1772 -3856 1824
rect -3844 1772 -3792 1824
rect -3592 1772 -3540 1824
rect -3528 1772 -3476 1824
rect -3276 1772 -3224 1824
rect -3212 1772 -3160 1824
rect -2960 1772 -2908 1824
rect -2896 1772 -2844 1824
rect -2644 1772 -2592 1824
rect -2580 1772 -2528 1824
rect -2328 1772 -2276 1824
rect -2264 1772 -2212 1824
rect -2012 1772 -1960 1824
rect -1948 1772 -1896 1824
rect -1696 1772 -1644 1824
rect -1632 1772 -1580 1824
rect -1380 1772 -1328 1824
rect -1316 1772 -1264 1824
rect -1064 1772 -1012 1824
rect -1000 1772 -948 1824
rect -748 1772 -696 1824
rect -684 1772 -632 1824
rect -432 1772 -380 1824
rect -368 1772 -316 1824
rect -116 1772 -64 1824
rect -52 1772 0 1824
rect 200 1772 252 1824
rect 264 1772 316 1824
rect 516 1772 568 1824
rect 580 1772 632 1824
rect 832 1772 884 1824
rect 896 1772 948 1824
rect 1148 1772 1200 1824
rect 1212 1772 1264 1824
rect 1464 1772 1516 1824
rect 1528 1772 1580 1824
rect 1780 1772 1832 1824
rect 1844 1772 1896 1824
rect 2096 1772 2148 1824
rect 2160 1772 2212 1824
rect -4036 1399 -3856 1400
rect -4036 1221 -4035 1399
rect -4035 1221 -3857 1399
rect -3857 1221 -3856 1399
rect -4036 1220 -3856 1221
rect -4343 932 -4342 1176
rect -4342 932 -4164 1176
rect -4164 932 -4163 1176
rect -4098 599 -3854 779
rect 2550 1508 2666 6104
rect -3173 1366 1295 1401
rect -3173 1260 1295 1366
rect -3173 1221 1295 1260
rect -3672 437 -3620 489
rect -3608 437 -3556 489
rect -2507 437 -2455 489
rect -2443 437 -2391 489
rect -2379 437 -2327 489
rect -2315 437 -2263 489
rect -2251 437 -2199 489
rect -2187 437 -2135 489
rect -3210 227 -3158 279
rect -3146 227 -3094 279
rect -3828 161 -3776 213
rect -3828 97 -3776 149
rect -4344 -307 -4164 1
rect -3861 -465 -3809 -413
rect -3797 -465 -3745 -413
rect -3214 -122 -3162 -70
rect -3214 -186 -3162 -134
rect -3214 -250 -3162 -198
rect -1338 435 -1286 487
rect -1274 435 -1222 487
rect -1210 435 -1158 487
rect -1146 435 -1094 487
rect -1082 435 -1030 487
rect -1018 435 -966 487
rect -2777 323 -2725 375
rect -2713 323 -2661 375
rect -2776 -122 -2724 -70
rect -2776 -186 -2724 -134
rect -2776 -250 -2724 -198
rect -1909 227 -1857 279
rect -1845 227 -1793 279
rect -2264 28 -2212 80
rect -2178 -119 -2126 -67
rect -2178 -183 -2126 -131
rect -2178 -247 -2126 -195
rect -1907 -120 -1855 -68
rect -1907 -184 -1855 -132
rect -1907 -248 -1855 -196
rect -1477 323 -1425 375
rect -1413 323 -1361 375
rect -1478 -119 -1426 -67
rect -1478 -183 -1426 -131
rect -1478 -247 -1426 -195
rect -592 780 -540 832
rect -592 716 -540 768
rect -592 652 -540 704
rect -654 323 -602 375
rect -590 323 -538 375
rect -526 323 -474 375
rect -961 28 -909 80
rect -7 778 45 830
rect -7 714 45 766
rect -7 650 45 702
rect -75 227 -23 279
rect -11 227 41 279
rect 53 227 105 279
rect 415 778 467 830
rect 415 714 467 766
rect 415 650 467 702
rect 735 781 787 833
rect 735 717 787 769
rect 735 653 787 705
rect 1003 746 1055 798
rect 1003 682 1055 734
rect -874 -119 -822 -67
rect -874 -183 -822 -131
rect -874 -247 -822 -195
rect -694 -465 -642 -413
rect -630 -465 -578 -413
rect 257 -164 309 -112
rect 257 -228 309 -176
rect 415 -144 467 -92
rect 415 -208 467 -156
rect 576 -162 628 -110
rect 576 -226 628 -174
rect 732 -144 784 -92
rect 732 -208 784 -156
rect 894 -161 946 -109
rect 894 -225 946 -173
rect 1045 -161 1097 -109
rect 1045 -225 1097 -173
rect 1755 435 1807 487
rect 1819 435 1871 487
rect 1883 435 1935 487
rect 2147 1401 2327 1402
rect 2147 1223 2148 1401
rect 2148 1223 2326 1401
rect 2326 1223 2327 1401
rect 2147 1222 2327 1223
rect 1599 122 1651 174
rect 1663 122 1715 174
rect 1467 7 1519 59
rect 1467 -57 1519 -5
rect 1327 -159 1379 -107
rect 1327 -223 1379 -171
rect 1467 -121 1519 -69
rect 1467 -185 1519 -133
rect 1467 -249 1519 -197
rect 1467 -313 1519 -261
rect 2550 694 2666 1002
rect 2478 408 2658 588
rect 2478 -82 2658 98
rect -3657 -583 -3605 -574
rect -3657 -617 -3652 -583
rect -3652 -617 -3618 -583
rect -3618 -617 -3605 -583
rect -3657 -626 -3605 -617
rect -3593 -583 -3541 -574
rect -3593 -617 -3580 -583
rect -3580 -617 -3546 -583
rect -3546 -617 -3541 -583
rect -3593 -626 -3541 -617
rect -3529 -583 -3477 -574
rect -3465 -583 -3413 -574
rect -3401 -583 -3349 -574
rect -3337 -583 -3285 -574
rect -3273 -583 -3221 -574
rect -3209 -583 -3157 -574
rect -3145 -583 -3093 -574
rect -3529 -617 -3508 -583
rect -3508 -617 -3477 -583
rect -3465 -617 -3436 -583
rect -3436 -617 -3413 -583
rect -3401 -617 -3364 -583
rect -3364 -617 -3349 -583
rect -3337 -617 -3330 -583
rect -3330 -617 -3292 -583
rect -3292 -617 -3285 -583
rect -3273 -617 -3258 -583
rect -3258 -617 -3221 -583
rect -3209 -617 -3186 -583
rect -3186 -617 -3157 -583
rect -3145 -617 -3114 -583
rect -3114 -617 -3093 -583
rect -3529 -626 -3477 -617
rect -3465 -626 -3413 -617
rect -3401 -626 -3349 -617
rect -3337 -626 -3285 -617
rect -3273 -626 -3221 -617
rect -3209 -626 -3157 -617
rect -3145 -626 -3093 -617
rect -3081 -583 -3029 -574
rect -3081 -617 -3076 -583
rect -3076 -617 -3042 -583
rect -3042 -617 -3029 -583
rect -3081 -626 -3029 -617
rect -3017 -583 -2965 -574
rect -3017 -617 -3004 -583
rect -3004 -617 -2970 -583
rect -2970 -617 -2965 -583
rect -3017 -626 -2965 -617
rect -2953 -583 -2901 -574
rect -2889 -583 -2837 -574
rect -2825 -583 -2773 -574
rect -2761 -583 -2709 -574
rect -2697 -583 -2645 -574
rect -2633 -583 -2581 -574
rect -2569 -583 -2517 -574
rect -2953 -617 -2932 -583
rect -2932 -617 -2901 -583
rect -2889 -617 -2860 -583
rect -2860 -617 -2837 -583
rect -2825 -617 -2788 -583
rect -2788 -617 -2773 -583
rect -2761 -617 -2754 -583
rect -2754 -617 -2716 -583
rect -2716 -617 -2709 -583
rect -2697 -617 -2682 -583
rect -2682 -617 -2645 -583
rect -2633 -617 -2610 -583
rect -2610 -617 -2581 -583
rect -2569 -617 -2538 -583
rect -2538 -617 -2517 -583
rect -2953 -626 -2901 -617
rect -2889 -626 -2837 -617
rect -2825 -626 -2773 -617
rect -2761 -626 -2709 -617
rect -2697 -626 -2645 -617
rect -2633 -626 -2581 -617
rect -2569 -626 -2517 -617
rect -2505 -583 -2453 -574
rect -2505 -617 -2500 -583
rect -2500 -617 -2466 -583
rect -2466 -617 -2453 -583
rect -2505 -626 -2453 -617
rect -2441 -583 -2389 -574
rect -2441 -617 -2428 -583
rect -2428 -617 -2394 -583
rect -2394 -617 -2389 -583
rect -2441 -626 -2389 -617
rect -2377 -583 -2325 -574
rect -2313 -583 -2261 -574
rect -2249 -583 -2197 -574
rect -2185 -583 -2133 -574
rect -2121 -583 -2069 -574
rect -2057 -583 -2005 -574
rect -1993 -583 -1941 -574
rect -2377 -617 -2356 -583
rect -2356 -617 -2325 -583
rect -2313 -617 -2284 -583
rect -2284 -617 -2261 -583
rect -2249 -617 -2212 -583
rect -2212 -617 -2197 -583
rect -2185 -617 -2178 -583
rect -2178 -617 -2140 -583
rect -2140 -617 -2133 -583
rect -2121 -617 -2106 -583
rect -2106 -617 -2069 -583
rect -2057 -617 -2034 -583
rect -2034 -617 -2005 -583
rect -1993 -617 -1962 -583
rect -1962 -617 -1941 -583
rect -2377 -626 -2325 -617
rect -2313 -626 -2261 -617
rect -2249 -626 -2197 -617
rect -2185 -626 -2133 -617
rect -2121 -626 -2069 -617
rect -2057 -626 -2005 -617
rect -1993 -626 -1941 -617
rect -1929 -583 -1877 -574
rect -1929 -617 -1924 -583
rect -1924 -617 -1890 -583
rect -1890 -617 -1877 -583
rect -1929 -626 -1877 -617
rect -1865 -583 -1813 -574
rect -1865 -617 -1852 -583
rect -1852 -617 -1818 -583
rect -1818 -617 -1813 -583
rect -1865 -626 -1813 -617
rect -1801 -583 -1749 -574
rect -1737 -583 -1685 -574
rect -1673 -583 -1621 -574
rect -1609 -583 -1557 -574
rect -1545 -583 -1493 -574
rect -1481 -583 -1429 -574
rect -1417 -583 -1365 -574
rect -1801 -617 -1780 -583
rect -1780 -617 -1749 -583
rect -1737 -617 -1708 -583
rect -1708 -617 -1685 -583
rect -1673 -617 -1636 -583
rect -1636 -617 -1621 -583
rect -1609 -617 -1602 -583
rect -1602 -617 -1564 -583
rect -1564 -617 -1557 -583
rect -1545 -617 -1530 -583
rect -1530 -617 -1493 -583
rect -1481 -617 -1458 -583
rect -1458 -617 -1429 -583
rect -1417 -617 -1386 -583
rect -1386 -617 -1365 -583
rect -1801 -626 -1749 -617
rect -1737 -626 -1685 -617
rect -1673 -626 -1621 -617
rect -1609 -626 -1557 -617
rect -1545 -626 -1493 -617
rect -1481 -626 -1429 -617
rect -1417 -626 -1365 -617
rect -1353 -583 -1301 -574
rect -1353 -617 -1348 -583
rect -1348 -617 -1314 -583
rect -1314 -617 -1301 -583
rect -1353 -626 -1301 -617
rect -1289 -583 -1237 -574
rect -1289 -617 -1276 -583
rect -1276 -617 -1242 -583
rect -1242 -617 -1237 -583
rect -1289 -626 -1237 -617
rect -1225 -583 -1173 -574
rect -1161 -583 -1109 -574
rect -1097 -583 -1045 -574
rect -1033 -583 -981 -574
rect -969 -583 -917 -574
rect -905 -583 -853 -574
rect -841 -583 -789 -574
rect -1225 -617 -1204 -583
rect -1204 -617 -1173 -583
rect -1161 -617 -1132 -583
rect -1132 -617 -1109 -583
rect -1097 -617 -1060 -583
rect -1060 -617 -1045 -583
rect -1033 -617 -1026 -583
rect -1026 -617 -988 -583
rect -988 -617 -981 -583
rect -969 -617 -954 -583
rect -954 -617 -917 -583
rect -905 -617 -882 -583
rect -882 -617 -853 -583
rect -841 -617 -810 -583
rect -810 -617 -789 -583
rect -1225 -626 -1173 -617
rect -1161 -626 -1109 -617
rect -1097 -626 -1045 -617
rect -1033 -626 -981 -617
rect -969 -626 -917 -617
rect -905 -626 -853 -617
rect -841 -626 -789 -617
rect -777 -583 -725 -574
rect -777 -617 -772 -583
rect -772 -617 -738 -583
rect -738 -617 -725 -583
rect -777 -626 -725 -617
rect -713 -583 -661 -574
rect -713 -617 -700 -583
rect -700 -617 -666 -583
rect -666 -617 -661 -583
rect -713 -626 -661 -617
rect -649 -583 -597 -574
rect -585 -583 -533 -574
rect -521 -583 -469 -574
rect -457 -583 -405 -574
rect -393 -583 -341 -574
rect -329 -583 -277 -574
rect -265 -583 -213 -574
rect -649 -617 -628 -583
rect -628 -617 -597 -583
rect -585 -617 -556 -583
rect -556 -617 -533 -583
rect -521 -617 -484 -583
rect -484 -617 -469 -583
rect -457 -617 -450 -583
rect -450 -617 -412 -583
rect -412 -617 -405 -583
rect -393 -617 -378 -583
rect -378 -617 -341 -583
rect -329 -617 -306 -583
rect -306 -617 -277 -583
rect -265 -617 -234 -583
rect -234 -617 -213 -583
rect -649 -626 -597 -617
rect -585 -626 -533 -617
rect -521 -626 -469 -617
rect -457 -626 -405 -617
rect -393 -626 -341 -617
rect -329 -626 -277 -617
rect -265 -626 -213 -617
rect -201 -583 -149 -574
rect -201 -617 -196 -583
rect -196 -617 -162 -583
rect -162 -617 -149 -583
rect -201 -626 -149 -617
rect -137 -583 -85 -574
rect -137 -617 -124 -583
rect -124 -617 -90 -583
rect -90 -617 -85 -583
rect -137 -626 -85 -617
rect -73 -583 -21 -574
rect -9 -583 43 -574
rect 55 -583 107 -574
rect 119 -583 171 -574
rect 183 -583 235 -574
rect 247 -583 299 -574
rect 311 -583 363 -574
rect -73 -617 -52 -583
rect -52 -617 -21 -583
rect -9 -617 20 -583
rect 20 -617 43 -583
rect 55 -617 92 -583
rect 92 -617 107 -583
rect 119 -617 126 -583
rect 126 -617 164 -583
rect 164 -617 171 -583
rect 183 -617 198 -583
rect 198 -617 235 -583
rect 247 -617 270 -583
rect 270 -617 299 -583
rect 311 -617 342 -583
rect 342 -617 363 -583
rect -73 -626 -21 -617
rect -9 -626 43 -617
rect 55 -626 107 -617
rect 119 -626 171 -617
rect 183 -626 235 -617
rect 247 -626 299 -617
rect 311 -626 363 -617
rect 375 -583 427 -574
rect 375 -617 380 -583
rect 380 -617 414 -583
rect 414 -617 427 -583
rect 375 -626 427 -617
rect 439 -583 491 -574
rect 439 -617 452 -583
rect 452 -617 486 -583
rect 486 -617 491 -583
rect 439 -626 491 -617
rect 503 -583 555 -574
rect 567 -583 619 -574
rect 631 -583 683 -574
rect 695 -583 747 -574
rect 759 -583 811 -574
rect 823 -583 875 -574
rect 887 -583 939 -574
rect 503 -617 524 -583
rect 524 -617 555 -583
rect 567 -617 596 -583
rect 596 -617 619 -583
rect 631 -617 668 -583
rect 668 -617 683 -583
rect 695 -617 702 -583
rect 702 -617 740 -583
rect 740 -617 747 -583
rect 759 -617 774 -583
rect 774 -617 811 -583
rect 823 -617 846 -583
rect 846 -617 875 -583
rect 887 -617 918 -583
rect 918 -617 939 -583
rect 503 -626 555 -617
rect 567 -626 619 -617
rect 631 -626 683 -617
rect 695 -626 747 -617
rect 759 -626 811 -617
rect 823 -626 875 -617
rect 887 -626 939 -617
rect 951 -583 1003 -574
rect 951 -617 956 -583
rect 956 -617 990 -583
rect 990 -617 1003 -583
rect 951 -626 1003 -617
rect 1015 -583 1067 -574
rect 1015 -617 1028 -583
rect 1028 -617 1062 -583
rect 1062 -617 1067 -583
rect 1015 -626 1067 -617
rect 1079 -583 1131 -574
rect 1143 -583 1195 -574
rect 1207 -583 1259 -574
rect 1271 -583 1323 -574
rect 1335 -583 1387 -574
rect 1399 -583 1451 -574
rect 1463 -583 1515 -574
rect 1079 -617 1100 -583
rect 1100 -617 1131 -583
rect 1143 -617 1172 -583
rect 1172 -617 1195 -583
rect 1207 -617 1244 -583
rect 1244 -617 1259 -583
rect 1271 -617 1278 -583
rect 1278 -617 1316 -583
rect 1316 -617 1323 -583
rect 1335 -617 1350 -583
rect 1350 -617 1387 -583
rect 1399 -617 1422 -583
rect 1422 -617 1451 -583
rect 1463 -617 1494 -583
rect 1494 -617 1515 -583
rect 1079 -626 1131 -617
rect 1143 -626 1195 -617
rect 1207 -626 1259 -617
rect 1271 -626 1323 -617
rect 1335 -626 1387 -617
rect 1399 -626 1451 -617
rect 1463 -626 1515 -617
rect 1527 -583 1579 -574
rect 1527 -617 1532 -583
rect 1532 -617 1566 -583
rect 1566 -617 1579 -583
rect 1527 -626 1579 -617
rect 1591 -583 1643 -574
rect 1591 -617 1604 -583
rect 1604 -617 1638 -583
rect 1638 -617 1643 -583
rect 1591 -626 1643 -617
rect 1655 -583 1707 -574
rect 1719 -583 1771 -574
rect 1783 -583 1835 -574
rect 1847 -583 1899 -574
rect 1911 -583 1963 -574
rect 1975 -583 2027 -574
rect 2039 -583 2091 -574
rect 1655 -617 1676 -583
rect 1676 -617 1707 -583
rect 1719 -617 1748 -583
rect 1748 -617 1771 -583
rect 1783 -617 1820 -583
rect 1820 -617 1835 -583
rect 1847 -617 1854 -583
rect 1854 -617 1892 -583
rect 1892 -617 1899 -583
rect 1911 -617 1926 -583
rect 1926 -617 1963 -583
rect 1975 -617 1998 -583
rect 1998 -617 2027 -583
rect 2039 -617 2070 -583
rect 2070 -617 2091 -583
rect 1655 -626 1707 -617
rect 1719 -626 1771 -617
rect 1783 -626 1835 -617
rect 1847 -626 1899 -617
rect 1911 -626 1963 -617
rect 1975 -626 2027 -617
rect 2039 -626 2091 -617
rect 2103 -583 2155 -574
rect 2103 -617 2108 -583
rect 2108 -617 2142 -583
rect 2142 -617 2155 -583
rect 2103 -626 2155 -617
rect 2167 -583 2219 -574
rect 2167 -617 2180 -583
rect 2180 -617 2214 -583
rect 2214 -617 2219 -583
rect 2167 -626 2219 -617
rect -4066 -936 -4014 -884
rect -4002 -936 -3950 -884
rect -3750 -936 -3698 -884
rect -3686 -936 -3634 -884
rect -3434 -936 -3382 -884
rect -3370 -936 -3318 -884
rect -3118 -936 -3066 -884
rect -3054 -936 -3002 -884
rect -2802 -936 -2750 -884
rect -2738 -936 -2686 -884
rect -2486 -936 -2434 -884
rect -2422 -936 -2370 -884
rect -2170 -936 -2118 -884
rect -2106 -936 -2054 -884
rect -1854 -936 -1802 -884
rect -1790 -936 -1738 -884
rect -1538 -936 -1486 -884
rect -1474 -936 -1422 -884
rect -1222 -936 -1170 -884
rect -1158 -936 -1106 -884
rect -906 -936 -854 -884
rect -842 -936 -790 -884
rect -590 -936 -538 -884
rect -526 -936 -474 -884
rect -274 -936 -222 -884
rect -210 -936 -158 -884
rect 42 -936 94 -884
rect 106 -936 158 -884
rect 358 -936 410 -884
rect 422 -936 474 -884
rect 674 -936 726 -884
rect 738 -936 790 -884
rect 990 -936 1042 -884
rect 1054 -936 1106 -884
rect 1306 -936 1358 -884
rect 1370 -936 1422 -884
rect 1622 -936 1674 -884
rect 1686 -936 1738 -884
rect 1938 -936 1990 -884
rect 2002 -936 2054 -884
rect 2254 -936 2306 -884
rect 2318 -936 2370 -884
rect -3908 -1061 -3856 -1009
rect -3844 -1061 -3792 -1009
rect -3592 -1061 -3540 -1009
rect -3528 -1061 -3476 -1009
rect -3276 -1061 -3224 -1009
rect -3212 -1061 -3160 -1009
rect -2960 -1061 -2908 -1009
rect -2896 -1061 -2844 -1009
rect -2644 -1061 -2592 -1009
rect -2580 -1061 -2528 -1009
rect -2328 -1061 -2276 -1009
rect -2264 -1061 -2212 -1009
rect -2012 -1061 -1960 -1009
rect -1948 -1061 -1896 -1009
rect -1696 -1061 -1644 -1009
rect -1632 -1061 -1580 -1009
rect -1380 -1061 -1328 -1009
rect -1316 -1061 -1264 -1009
rect -1064 -1061 -1012 -1009
rect -1000 -1061 -948 -1009
rect -748 -1061 -696 -1009
rect -684 -1061 -632 -1009
rect -432 -1061 -380 -1009
rect -368 -1061 -316 -1009
rect -116 -1061 -64 -1009
rect -52 -1061 0 -1009
rect 200 -1061 252 -1009
rect 264 -1061 316 -1009
rect 516 -1061 568 -1009
rect 580 -1061 632 -1009
rect 832 -1061 884 -1009
rect 896 -1061 948 -1009
rect 1148 -1061 1200 -1009
rect 1212 -1061 1264 -1009
rect 1464 -1061 1516 -1009
rect 1528 -1061 1580 -1009
rect 1780 -1061 1832 -1009
rect 1844 -1061 1896 -1009
rect 2096 -1061 2148 -1009
rect 2160 -1061 2212 -1009
rect -4066 -1354 -4014 -1302
rect -4002 -1354 -3950 -1302
rect -3750 -1354 -3698 -1302
rect -3686 -1354 -3634 -1302
rect -3434 -1354 -3382 -1302
rect -3370 -1354 -3318 -1302
rect -3118 -1354 -3066 -1302
rect -3054 -1354 -3002 -1302
rect -2802 -1354 -2750 -1302
rect -2738 -1354 -2686 -1302
rect -2486 -1354 -2434 -1302
rect -2422 -1354 -2370 -1302
rect -2170 -1354 -2118 -1302
rect -2106 -1354 -2054 -1302
rect -1854 -1354 -1802 -1302
rect -1790 -1354 -1738 -1302
rect -1538 -1354 -1486 -1302
rect -1474 -1354 -1422 -1302
rect -1222 -1354 -1170 -1302
rect -1158 -1354 -1106 -1302
rect -906 -1354 -854 -1302
rect -842 -1354 -790 -1302
rect -590 -1354 -538 -1302
rect -526 -1354 -474 -1302
rect -274 -1354 -222 -1302
rect -210 -1354 -158 -1302
rect 42 -1354 94 -1302
rect 106 -1354 158 -1302
rect 358 -1354 410 -1302
rect 422 -1354 474 -1302
rect 674 -1354 726 -1302
rect 738 -1354 790 -1302
rect 990 -1354 1042 -1302
rect 1054 -1354 1106 -1302
rect 1306 -1354 1358 -1302
rect 1370 -1354 1422 -1302
rect 1622 -1354 1674 -1302
rect 1686 -1354 1738 -1302
rect 1938 -1354 1990 -1302
rect 2002 -1354 2054 -1302
rect 2254 -1354 2306 -1302
rect 2318 -1354 2370 -1302
rect -3908 -1479 -3856 -1427
rect -3844 -1479 -3792 -1427
rect -3592 -1479 -3540 -1427
rect -3528 -1479 -3476 -1427
rect -3276 -1479 -3224 -1427
rect -3212 -1479 -3160 -1427
rect -2960 -1479 -2908 -1427
rect -2896 -1479 -2844 -1427
rect -2644 -1479 -2592 -1427
rect -2580 -1479 -2528 -1427
rect -2328 -1479 -2276 -1427
rect -2264 -1479 -2212 -1427
rect -2012 -1479 -1960 -1427
rect -1948 -1479 -1896 -1427
rect -1696 -1479 -1644 -1427
rect -1632 -1479 -1580 -1427
rect -1380 -1479 -1328 -1427
rect -1316 -1479 -1264 -1427
rect -1064 -1479 -1012 -1427
rect -1000 -1479 -948 -1427
rect -748 -1479 -696 -1427
rect -684 -1479 -632 -1427
rect -432 -1479 -380 -1427
rect -368 -1479 -316 -1427
rect -116 -1479 -64 -1427
rect -52 -1479 0 -1427
rect 200 -1479 252 -1427
rect 264 -1479 316 -1427
rect 516 -1479 568 -1427
rect 580 -1479 632 -1427
rect 832 -1479 884 -1427
rect 896 -1479 948 -1427
rect 1148 -1479 1200 -1427
rect 1212 -1479 1264 -1427
rect 1464 -1479 1516 -1427
rect 1528 -1479 1580 -1427
rect 1780 -1479 1832 -1427
rect 1844 -1479 1896 -1427
rect 2096 -1479 2148 -1427
rect 2160 -1479 2212 -1427
rect -4066 -1772 -4014 -1720
rect -4002 -1772 -3950 -1720
rect -3750 -1772 -3698 -1720
rect -3686 -1772 -3634 -1720
rect -3434 -1772 -3382 -1720
rect -3370 -1772 -3318 -1720
rect -3118 -1772 -3066 -1720
rect -3054 -1772 -3002 -1720
rect -2802 -1772 -2750 -1720
rect -2738 -1772 -2686 -1720
rect -2486 -1772 -2434 -1720
rect -2422 -1772 -2370 -1720
rect -2170 -1772 -2118 -1720
rect -2106 -1772 -2054 -1720
rect -1854 -1772 -1802 -1720
rect -1790 -1772 -1738 -1720
rect -1538 -1772 -1486 -1720
rect -1474 -1772 -1422 -1720
rect -1222 -1772 -1170 -1720
rect -1158 -1772 -1106 -1720
rect -906 -1772 -854 -1720
rect -842 -1772 -790 -1720
rect -590 -1772 -538 -1720
rect -526 -1772 -474 -1720
rect -274 -1772 -222 -1720
rect -210 -1772 -158 -1720
rect 42 -1772 94 -1720
rect 106 -1772 158 -1720
rect 358 -1772 410 -1720
rect 422 -1772 474 -1720
rect 674 -1772 726 -1720
rect 738 -1772 790 -1720
rect 990 -1772 1042 -1720
rect 1054 -1772 1106 -1720
rect 1306 -1772 1358 -1720
rect 1370 -1772 1422 -1720
rect 1622 -1772 1674 -1720
rect 1686 -1772 1738 -1720
rect 1938 -1772 1990 -1720
rect 2002 -1772 2054 -1720
rect 2254 -1772 2306 -1720
rect 2318 -1772 2370 -1720
rect -3908 -1897 -3856 -1845
rect -3844 -1897 -3792 -1845
rect -3592 -1897 -3540 -1845
rect -3528 -1897 -3476 -1845
rect -3276 -1897 -3224 -1845
rect -3212 -1897 -3160 -1845
rect -2960 -1897 -2908 -1845
rect -2896 -1897 -2844 -1845
rect -2644 -1897 -2592 -1845
rect -2580 -1897 -2528 -1845
rect -2328 -1897 -2276 -1845
rect -2264 -1897 -2212 -1845
rect -2012 -1897 -1960 -1845
rect -1948 -1897 -1896 -1845
rect -1696 -1897 -1644 -1845
rect -1632 -1897 -1580 -1845
rect -1380 -1897 -1328 -1845
rect -1316 -1897 -1264 -1845
rect -1064 -1897 -1012 -1845
rect -1000 -1897 -948 -1845
rect -748 -1897 -696 -1845
rect -684 -1897 -632 -1845
rect -432 -1897 -380 -1845
rect -368 -1897 -316 -1845
rect -116 -1897 -64 -1845
rect -52 -1897 0 -1845
rect 200 -1897 252 -1845
rect 264 -1897 316 -1845
rect 516 -1897 568 -1845
rect 580 -1897 632 -1845
rect 832 -1897 884 -1845
rect 896 -1897 948 -1845
rect 1148 -1897 1200 -1845
rect 1212 -1897 1264 -1845
rect 1464 -1897 1516 -1845
rect 1528 -1897 1580 -1845
rect 1780 -1897 1832 -1845
rect 1844 -1897 1896 -1845
rect 2096 -1897 2148 -1845
rect 2160 -1897 2212 -1845
rect -4380 -2439 -4136 -2131
rect 1631 -3412 2195 -3296
rect 2638 -3286 2682 -3234
rect 2682 -3286 2690 -3234
rect 2638 -3350 2682 -3298
rect 2682 -3350 2690 -3298
rect 2638 -3414 2682 -3362
rect 2682 -3414 2690 -3362
rect 2638 -3478 2682 -3426
rect 2682 -3478 2690 -3426
<< metal2 >>
rect -4362 6475 2685 6535
rect -4362 6359 -4326 6475
rect 2638 6359 2685 6475
rect -4362 6313 2685 6359
rect -4362 5931 -4140 6313
rect -4081 6104 2683 6130
rect -4081 6049 2550 6104
rect -4081 5997 -4066 6049
rect -4014 5997 -4002 6049
rect -3950 5997 -3750 6049
rect -3698 5997 -3686 6049
rect -3634 5997 -3434 6049
rect -3382 5997 -3370 6049
rect -3318 5997 -3118 6049
rect -3066 5997 -3054 6049
rect -3002 5997 -2802 6049
rect -2750 5997 -2738 6049
rect -2686 5997 -2486 6049
rect -2434 5997 -2422 6049
rect -2370 5997 -2170 6049
rect -2118 5997 -2106 6049
rect -2054 5997 -1854 6049
rect -1802 5997 -1790 6049
rect -1738 5997 -1538 6049
rect -1486 5997 -1474 6049
rect -1422 5997 -1222 6049
rect -1170 5997 -1158 6049
rect -1106 5997 -906 6049
rect -854 5997 -842 6049
rect -790 5997 -590 6049
rect -538 5997 -526 6049
rect -474 5997 -274 6049
rect -222 5997 -210 6049
rect -158 5997 42 6049
rect 94 5997 106 6049
rect 158 5997 358 6049
rect 410 5997 422 6049
rect 474 5997 674 6049
rect 726 5997 738 6049
rect 790 5997 990 6049
rect 1042 5997 1054 6049
rect 1106 5997 1306 6049
rect 1358 5997 1370 6049
rect 1422 5997 1622 6049
rect 1674 5997 1686 6049
rect 1738 5997 1938 6049
rect 1990 5997 2002 6049
rect 2054 5997 2254 6049
rect 2306 5997 2318 6049
rect 2370 5997 2550 6049
rect -4081 5991 2550 5997
rect -4362 5930 -4081 5931
rect -4362 5924 2399 5930
rect -4362 5872 -3908 5924
rect -3856 5872 -3844 5924
rect -3792 5872 -3592 5924
rect -3540 5872 -3528 5924
rect -3476 5872 -3276 5924
rect -3224 5872 -3212 5924
rect -3160 5872 -2960 5924
rect -2908 5872 -2896 5924
rect -2844 5872 -2644 5924
rect -2592 5872 -2580 5924
rect -2528 5872 -2328 5924
rect -2276 5872 -2264 5924
rect -2212 5872 -2012 5924
rect -1960 5872 -1948 5924
rect -1896 5872 -1696 5924
rect -1644 5872 -1632 5924
rect -1580 5872 -1380 5924
rect -1328 5872 -1316 5924
rect -1264 5872 -1064 5924
rect -1012 5872 -1000 5924
rect -948 5872 -748 5924
rect -696 5872 -684 5924
rect -632 5872 -432 5924
rect -380 5872 -368 5924
rect -316 5872 -116 5924
rect -64 5872 -52 5924
rect 0 5872 200 5924
rect 252 5872 264 5924
rect 316 5872 516 5924
rect 568 5872 580 5924
rect 632 5872 832 5924
rect 884 5872 896 5924
rect 948 5872 1148 5924
rect 1200 5872 1212 5924
rect 1264 5872 1464 5924
rect 1516 5872 1528 5924
rect 1580 5872 1780 5924
rect 1832 5872 1844 5924
rect 1896 5872 2096 5924
rect 2148 5872 2160 5924
rect 2212 5872 2399 5924
rect -4362 5792 2399 5872
rect -4362 5490 -4140 5792
rect -4081 5791 2399 5792
rect 2453 5690 2550 5991
rect -4081 5609 2550 5690
rect -4081 5557 -4066 5609
rect -4014 5557 -4002 5609
rect -3950 5557 -3750 5609
rect -3698 5557 -3686 5609
rect -3634 5557 -3434 5609
rect -3382 5557 -3370 5609
rect -3318 5557 -3118 5609
rect -3066 5557 -3054 5609
rect -3002 5557 -2802 5609
rect -2750 5557 -2738 5609
rect -2686 5557 -2486 5609
rect -2434 5557 -2422 5609
rect -2370 5557 -2170 5609
rect -2118 5557 -2106 5609
rect -2054 5557 -1854 5609
rect -1802 5557 -1790 5609
rect -1738 5557 -1538 5609
rect -1486 5557 -1474 5609
rect -1422 5557 -1222 5609
rect -1170 5557 -1158 5609
rect -1106 5557 -906 5609
rect -854 5557 -842 5609
rect -790 5557 -590 5609
rect -538 5557 -526 5609
rect -474 5557 -274 5609
rect -222 5557 -210 5609
rect -158 5557 42 5609
rect 94 5557 106 5609
rect 158 5557 358 5609
rect 410 5557 422 5609
rect 474 5557 674 5609
rect 726 5557 738 5609
rect 790 5557 990 5609
rect 1042 5557 1054 5609
rect 1106 5557 1306 5609
rect 1358 5557 1370 5609
rect 1422 5557 1622 5609
rect 1674 5557 1686 5609
rect 1738 5557 1938 5609
rect 1990 5557 2002 5609
rect 2054 5557 2254 5609
rect 2306 5557 2318 5609
rect 2370 5557 2550 5609
rect -4081 5551 2550 5557
rect -4362 5484 2399 5490
rect -4362 5432 -3908 5484
rect -3856 5432 -3844 5484
rect -3792 5432 -3592 5484
rect -3540 5432 -3528 5484
rect -3476 5432 -3276 5484
rect -3224 5432 -3212 5484
rect -3160 5432 -2960 5484
rect -2908 5432 -2896 5484
rect -2844 5432 -2644 5484
rect -2592 5432 -2580 5484
rect -2528 5432 -2328 5484
rect -2276 5432 -2264 5484
rect -2212 5432 -2012 5484
rect -1960 5432 -1948 5484
rect -1896 5432 -1696 5484
rect -1644 5432 -1632 5484
rect -1580 5432 -1380 5484
rect -1328 5432 -1316 5484
rect -1264 5432 -1064 5484
rect -1012 5432 -1000 5484
rect -948 5432 -748 5484
rect -696 5432 -684 5484
rect -632 5432 -432 5484
rect -380 5432 -368 5484
rect -316 5432 -116 5484
rect -64 5432 -52 5484
rect 0 5432 200 5484
rect 252 5432 264 5484
rect 316 5432 516 5484
rect 568 5432 580 5484
rect 632 5432 832 5484
rect 884 5432 896 5484
rect 948 5432 1148 5484
rect 1200 5432 1212 5484
rect 1264 5432 1464 5484
rect 1516 5432 1528 5484
rect 1580 5432 1780 5484
rect 1832 5432 1844 5484
rect 1896 5432 2096 5484
rect 2148 5432 2160 5484
rect 2212 5432 2399 5484
rect -4362 5351 2399 5432
rect -4362 5050 -4140 5351
rect 2453 5250 2550 5551
rect -4081 5169 2550 5250
rect -4081 5117 -4066 5169
rect -4014 5117 -4002 5169
rect -3950 5117 -3750 5169
rect -3698 5117 -3686 5169
rect -3634 5117 -3434 5169
rect -3382 5117 -3370 5169
rect -3318 5117 -3118 5169
rect -3066 5117 -3054 5169
rect -3002 5117 -2802 5169
rect -2750 5117 -2738 5169
rect -2686 5117 -2486 5169
rect -2434 5117 -2422 5169
rect -2370 5117 -2170 5169
rect -2118 5117 -2106 5169
rect -2054 5117 -1854 5169
rect -1802 5117 -1790 5169
rect -1738 5117 -1538 5169
rect -1486 5117 -1474 5169
rect -1422 5117 -1222 5169
rect -1170 5117 -1158 5169
rect -1106 5117 -906 5169
rect -854 5117 -842 5169
rect -790 5117 -590 5169
rect -538 5117 -526 5169
rect -474 5117 -274 5169
rect -222 5117 -210 5169
rect -158 5117 42 5169
rect 94 5117 106 5169
rect 158 5117 358 5169
rect 410 5117 422 5169
rect 474 5117 674 5169
rect 726 5117 738 5169
rect 790 5117 990 5169
rect 1042 5117 1054 5169
rect 1106 5117 1306 5169
rect 1358 5117 1370 5169
rect 1422 5117 1622 5169
rect 1674 5117 1686 5169
rect 1738 5117 1938 5169
rect 1990 5117 2002 5169
rect 2054 5117 2254 5169
rect 2306 5117 2318 5169
rect 2370 5117 2550 5169
rect -4081 5111 2550 5117
rect -4362 5044 2399 5050
rect -4362 4992 -3908 5044
rect -3856 4992 -3844 5044
rect -3792 4992 -3592 5044
rect -3540 4992 -3528 5044
rect -3476 4992 -3276 5044
rect -3224 4992 -3212 5044
rect -3160 4992 -2960 5044
rect -2908 4992 -2896 5044
rect -2844 4992 -2644 5044
rect -2592 4992 -2580 5044
rect -2528 4992 -2328 5044
rect -2276 4992 -2264 5044
rect -2212 4992 -2012 5044
rect -1960 4992 -1948 5044
rect -1896 4992 -1696 5044
rect -1644 4992 -1632 5044
rect -1580 4992 -1380 5044
rect -1328 4992 -1316 5044
rect -1264 4992 -1064 5044
rect -1012 4992 -1000 5044
rect -948 4992 -748 5044
rect -696 4992 -684 5044
rect -632 4992 -432 5044
rect -380 4992 -368 5044
rect -316 4992 -116 5044
rect -64 4992 -52 5044
rect 0 4992 200 5044
rect 252 4992 264 5044
rect 316 4992 516 5044
rect 568 4992 580 5044
rect 632 4992 832 5044
rect 884 4992 896 5044
rect 948 4992 1148 5044
rect 1200 4992 1212 5044
rect 1264 4992 1464 5044
rect 1516 4992 1528 5044
rect 1580 4992 1780 5044
rect 1832 4992 1844 5044
rect 1896 4992 2096 5044
rect 2148 4992 2160 5044
rect 2212 4992 2399 5044
rect -4362 4911 2399 4992
rect -4362 4615 -4140 4911
rect 2453 4815 2550 5111
rect -4081 4734 2550 4815
rect -4081 4682 -4066 4734
rect -4014 4682 -4002 4734
rect -3950 4682 -3750 4734
rect -3698 4682 -3686 4734
rect -3634 4682 -3434 4734
rect -3382 4682 -3370 4734
rect -3318 4682 -3118 4734
rect -3066 4682 -3054 4734
rect -3002 4682 -2802 4734
rect -2750 4682 -2738 4734
rect -2686 4682 -2486 4734
rect -2434 4682 -2422 4734
rect -2370 4682 -2170 4734
rect -2118 4682 -2106 4734
rect -2054 4682 -1854 4734
rect -1802 4682 -1790 4734
rect -1738 4682 -1538 4734
rect -1486 4682 -1474 4734
rect -1422 4682 -1222 4734
rect -1170 4682 -1158 4734
rect -1106 4682 -906 4734
rect -854 4682 -842 4734
rect -790 4682 -590 4734
rect -538 4682 -526 4734
rect -474 4682 -274 4734
rect -222 4682 -210 4734
rect -158 4682 42 4734
rect 94 4682 106 4734
rect 158 4682 358 4734
rect 410 4682 422 4734
rect 474 4682 674 4734
rect 726 4682 738 4734
rect 790 4682 990 4734
rect 1042 4682 1054 4734
rect 1106 4682 1306 4734
rect 1358 4682 1370 4734
rect 1422 4682 1622 4734
rect 1674 4682 1686 4734
rect 1738 4682 1938 4734
rect 1990 4682 2002 4734
rect 2054 4682 2254 4734
rect 2306 4682 2318 4734
rect 2370 4682 2550 4734
rect -4081 4676 2550 4682
rect -4362 4609 2399 4615
rect -4362 4557 -3908 4609
rect -3856 4557 -3844 4609
rect -3792 4557 -3592 4609
rect -3540 4557 -3528 4609
rect -3476 4557 -3276 4609
rect -3224 4557 -3212 4609
rect -3160 4557 -2960 4609
rect -2908 4557 -2896 4609
rect -2844 4557 -2644 4609
rect -2592 4557 -2580 4609
rect -2528 4557 -2328 4609
rect -2276 4557 -2264 4609
rect -2212 4557 -2012 4609
rect -1960 4557 -1948 4609
rect -1896 4557 -1696 4609
rect -1644 4557 -1632 4609
rect -1580 4557 -1380 4609
rect -1328 4557 -1316 4609
rect -1264 4557 -1064 4609
rect -1012 4557 -1000 4609
rect -948 4557 -748 4609
rect -696 4557 -684 4609
rect -632 4557 -432 4609
rect -380 4557 -368 4609
rect -316 4557 -116 4609
rect -64 4557 -52 4609
rect 0 4557 200 4609
rect 252 4557 264 4609
rect 316 4557 516 4609
rect 568 4557 580 4609
rect 632 4557 832 4609
rect 884 4557 896 4609
rect 948 4557 1148 4609
rect 1200 4557 1212 4609
rect 1264 4557 1464 4609
rect 1516 4557 1528 4609
rect 1580 4557 1780 4609
rect 1832 4557 1844 4609
rect 1896 4557 2096 4609
rect 2148 4557 2160 4609
rect 2212 4557 2399 4609
rect -4362 4476 2399 4557
rect -4362 4190 -4140 4476
rect 2453 4390 2550 4676
rect -4081 4309 2550 4390
rect -4081 4257 -4066 4309
rect -4014 4257 -4002 4309
rect -3950 4257 -3750 4309
rect -3698 4257 -3686 4309
rect -3634 4257 -3434 4309
rect -3382 4257 -3370 4309
rect -3318 4257 -3118 4309
rect -3066 4257 -3054 4309
rect -3002 4257 -2802 4309
rect -2750 4257 -2738 4309
rect -2686 4257 -2486 4309
rect -2434 4257 -2422 4309
rect -2370 4257 -2170 4309
rect -2118 4257 -2106 4309
rect -2054 4257 -1854 4309
rect -1802 4257 -1790 4309
rect -1738 4257 -1538 4309
rect -1486 4257 -1474 4309
rect -1422 4257 -1222 4309
rect -1170 4257 -1158 4309
rect -1106 4257 -906 4309
rect -854 4257 -842 4309
rect -790 4257 -590 4309
rect -538 4257 -526 4309
rect -474 4257 -274 4309
rect -222 4257 -210 4309
rect -158 4257 42 4309
rect 94 4257 106 4309
rect 158 4257 358 4309
rect 410 4257 422 4309
rect 474 4257 674 4309
rect 726 4257 738 4309
rect 790 4257 990 4309
rect 1042 4257 1054 4309
rect 1106 4257 1306 4309
rect 1358 4257 1370 4309
rect 1422 4257 1622 4309
rect 1674 4257 1686 4309
rect 1738 4257 1938 4309
rect 1990 4257 2002 4309
rect 2054 4257 2254 4309
rect 2306 4257 2318 4309
rect 2370 4257 2550 4309
rect -4081 4251 2550 4257
rect -4362 4184 2399 4190
rect -4362 4132 -3908 4184
rect -3856 4132 -3844 4184
rect -3792 4132 -3592 4184
rect -3540 4132 -3528 4184
rect -3476 4132 -3276 4184
rect -3224 4132 -3212 4184
rect -3160 4132 -2960 4184
rect -2908 4132 -2896 4184
rect -2844 4132 -2644 4184
rect -2592 4132 -2580 4184
rect -2528 4132 -2328 4184
rect -2276 4132 -2264 4184
rect -2212 4132 -2012 4184
rect -1960 4132 -1948 4184
rect -1896 4132 -1696 4184
rect -1644 4132 -1632 4184
rect -1580 4132 -1380 4184
rect -1328 4132 -1316 4184
rect -1264 4132 -1064 4184
rect -1012 4132 -1000 4184
rect -948 4132 -748 4184
rect -696 4132 -684 4184
rect -632 4132 -432 4184
rect -380 4132 -368 4184
rect -316 4132 -116 4184
rect -64 4132 -52 4184
rect 0 4132 200 4184
rect 252 4132 264 4184
rect 316 4132 516 4184
rect 568 4132 580 4184
rect 632 4132 832 4184
rect 884 4132 896 4184
rect 948 4132 1148 4184
rect 1200 4132 1212 4184
rect 1264 4132 1464 4184
rect 1516 4132 1528 4184
rect 1580 4132 1780 4184
rect 1832 4132 1844 4184
rect 1896 4132 2096 4184
rect 2148 4132 2160 4184
rect 2212 4132 2399 4184
rect -4362 4051 2399 4132
rect -4362 3941 -4140 4051
rect 2453 4002 2550 4251
rect 2470 3974 2550 4002
rect -4362 3937 2376 3941
rect -4362 3885 -4110 3937
rect -4058 3885 -4046 3937
rect -3994 3885 -3982 3937
rect -3930 3885 -3918 3937
rect -3866 3885 -3854 3937
rect -3802 3885 -3790 3937
rect -3738 3885 -3726 3937
rect -3674 3885 -3662 3937
rect -3610 3885 -3598 3937
rect -3546 3885 -3534 3937
rect -3482 3885 -3470 3937
rect -3418 3885 -3406 3937
rect -3354 3885 -3342 3937
rect -3290 3885 -3278 3937
rect -3226 3885 -3214 3937
rect -3162 3885 -3150 3937
rect -3098 3885 -3086 3937
rect -3034 3885 -3022 3937
rect -2970 3885 -2958 3937
rect -2906 3885 -2894 3937
rect -2842 3885 -2830 3937
rect -2778 3885 -2766 3937
rect -2714 3885 -2702 3937
rect -2650 3885 -2638 3937
rect -2586 3885 -2574 3937
rect -2522 3885 -2510 3937
rect -2458 3885 -2446 3937
rect -2394 3885 -2382 3937
rect -2330 3885 -2318 3937
rect -2266 3885 -2254 3937
rect -2202 3885 -2190 3937
rect -2138 3885 -2126 3937
rect -2074 3885 -2062 3937
rect -2010 3885 -1998 3937
rect -1946 3885 -1934 3937
rect -1882 3885 -1870 3937
rect -1818 3885 -1806 3937
rect -1754 3885 -1742 3937
rect -1690 3885 -1678 3937
rect -1626 3885 -1614 3937
rect -1562 3885 -1550 3937
rect -1498 3885 -1486 3937
rect -1434 3885 -1422 3937
rect -1370 3885 -1358 3937
rect -1306 3885 -1294 3937
rect -1242 3885 -1230 3937
rect -1178 3885 -1166 3937
rect -1114 3885 -1102 3937
rect -1050 3885 -1038 3937
rect -986 3885 -974 3937
rect -922 3885 -910 3937
rect -858 3885 -846 3937
rect -794 3885 -782 3937
rect -730 3885 -718 3937
rect -666 3885 -654 3937
rect -602 3885 -590 3937
rect -538 3885 -526 3937
rect -474 3885 -462 3937
rect -410 3885 -398 3937
rect -346 3885 -334 3937
rect -282 3885 -270 3937
rect -218 3885 -206 3937
rect -154 3885 -142 3937
rect -90 3885 -78 3937
rect -26 3885 -14 3937
rect 38 3885 50 3937
rect 102 3885 114 3937
rect 166 3885 178 3937
rect 230 3885 242 3937
rect 294 3885 306 3937
rect 358 3885 370 3937
rect 422 3885 434 3937
rect 486 3885 498 3937
rect 550 3885 562 3937
rect 614 3885 626 3937
rect 678 3885 690 3937
rect 742 3885 754 3937
rect 806 3885 818 3937
rect 870 3885 882 3937
rect 934 3885 946 3937
rect 998 3885 1010 3937
rect 1062 3885 1074 3937
rect 1126 3885 1138 3937
rect 1190 3885 1202 3937
rect 1254 3885 1266 3937
rect 1318 3885 1330 3937
rect 1382 3885 1394 3937
rect 1446 3885 1458 3937
rect 1510 3885 1522 3937
rect 1574 3885 1586 3937
rect 1638 3885 1650 3937
rect 1702 3885 1714 3937
rect 1766 3885 1778 3937
rect 1830 3885 1842 3937
rect 1894 3885 1906 3937
rect 1958 3885 1970 3937
rect 2022 3885 2034 3937
rect 2086 3885 2098 3937
rect 2150 3885 2162 3937
rect 2214 3885 2226 3937
rect 2278 3885 2290 3937
rect 2342 3885 2376 3937
rect -4362 3881 2376 3885
rect -4362 3570 -4140 3881
rect 2453 3770 2550 3974
rect -4081 3689 2550 3770
rect -4081 3637 -4066 3689
rect -4014 3637 -4002 3689
rect -3950 3637 -3750 3689
rect -3698 3637 -3686 3689
rect -3634 3637 -3434 3689
rect -3382 3637 -3370 3689
rect -3318 3637 -3118 3689
rect -3066 3637 -3054 3689
rect -3002 3637 -2802 3689
rect -2750 3637 -2738 3689
rect -2686 3637 -2486 3689
rect -2434 3637 -2422 3689
rect -2370 3637 -2170 3689
rect -2118 3637 -2106 3689
rect -2054 3637 -1854 3689
rect -1802 3637 -1790 3689
rect -1738 3637 -1538 3689
rect -1486 3637 -1474 3689
rect -1422 3637 -1222 3689
rect -1170 3637 -1158 3689
rect -1106 3637 -906 3689
rect -854 3637 -842 3689
rect -790 3637 -590 3689
rect -538 3637 -526 3689
rect -474 3637 -274 3689
rect -222 3637 -210 3689
rect -158 3637 42 3689
rect 94 3637 106 3689
rect 158 3637 358 3689
rect 410 3637 422 3689
rect 474 3637 674 3689
rect 726 3637 738 3689
rect 790 3637 990 3689
rect 1042 3637 1054 3689
rect 1106 3637 1306 3689
rect 1358 3637 1370 3689
rect 1422 3637 1622 3689
rect 1674 3637 1686 3689
rect 1738 3637 1938 3689
rect 1990 3637 2002 3689
rect 2054 3637 2254 3689
rect 2306 3637 2318 3689
rect 2370 3637 2550 3689
rect -4081 3631 2550 3637
rect -4362 3564 2399 3570
rect -4362 3512 -3908 3564
rect -3856 3512 -3844 3564
rect -3792 3512 -3592 3564
rect -3540 3512 -3528 3564
rect -3476 3512 -3276 3564
rect -3224 3512 -3212 3564
rect -3160 3512 -2960 3564
rect -2908 3512 -2896 3564
rect -2844 3512 -2644 3564
rect -2592 3512 -2580 3564
rect -2528 3512 -2328 3564
rect -2276 3512 -2264 3564
rect -2212 3512 -2012 3564
rect -1960 3512 -1948 3564
rect -1896 3512 -1696 3564
rect -1644 3512 -1632 3564
rect -1580 3512 -1380 3564
rect -1328 3512 -1316 3564
rect -1264 3512 -1064 3564
rect -1012 3512 -1000 3564
rect -948 3512 -748 3564
rect -696 3512 -684 3564
rect -632 3512 -432 3564
rect -380 3512 -368 3564
rect -316 3512 -116 3564
rect -64 3512 -52 3564
rect 0 3512 200 3564
rect 252 3512 264 3564
rect 316 3512 516 3564
rect 568 3512 580 3564
rect 632 3512 832 3564
rect 884 3512 896 3564
rect 948 3512 1148 3564
rect 1200 3512 1212 3564
rect 1264 3512 1464 3564
rect 1516 3512 1528 3564
rect 1580 3512 1780 3564
rect 1832 3512 1844 3564
rect 1896 3512 2096 3564
rect 2148 3512 2160 3564
rect 2212 3512 2399 3564
rect -4362 3431 2399 3512
rect -4362 3135 -4140 3431
rect 2453 3335 2550 3631
rect -4081 3254 2550 3335
rect -4081 3202 -4066 3254
rect -4014 3202 -4002 3254
rect -3950 3202 -3750 3254
rect -3698 3202 -3686 3254
rect -3634 3202 -3434 3254
rect -3382 3202 -3370 3254
rect -3318 3202 -3118 3254
rect -3066 3202 -3054 3254
rect -3002 3202 -2802 3254
rect -2750 3202 -2738 3254
rect -2686 3202 -2486 3254
rect -2434 3202 -2422 3254
rect -2370 3202 -2170 3254
rect -2118 3202 -2106 3254
rect -2054 3202 -1854 3254
rect -1802 3202 -1790 3254
rect -1738 3202 -1538 3254
rect -1486 3202 -1474 3254
rect -1422 3202 -1222 3254
rect -1170 3202 -1158 3254
rect -1106 3202 -906 3254
rect -854 3202 -842 3254
rect -790 3202 -590 3254
rect -538 3202 -526 3254
rect -474 3202 -274 3254
rect -222 3202 -210 3254
rect -158 3202 42 3254
rect 94 3202 106 3254
rect 158 3202 358 3254
rect 410 3202 422 3254
rect 474 3202 674 3254
rect 726 3202 738 3254
rect 790 3202 990 3254
rect 1042 3202 1054 3254
rect 1106 3202 1306 3254
rect 1358 3202 1370 3254
rect 1422 3202 1622 3254
rect 1674 3202 1686 3254
rect 1738 3202 1938 3254
rect 1990 3202 2002 3254
rect 2054 3202 2254 3254
rect 2306 3202 2318 3254
rect 2370 3202 2550 3254
rect -4081 3196 2550 3202
rect -4362 3129 2399 3135
rect -4362 3077 -3908 3129
rect -3856 3077 -3844 3129
rect -3792 3077 -3592 3129
rect -3540 3077 -3528 3129
rect -3476 3077 -3276 3129
rect -3224 3077 -3212 3129
rect -3160 3077 -2960 3129
rect -2908 3077 -2896 3129
rect -2844 3077 -2644 3129
rect -2592 3077 -2580 3129
rect -2528 3077 -2328 3129
rect -2276 3077 -2264 3129
rect -2212 3077 -2012 3129
rect -1960 3077 -1948 3129
rect -1896 3077 -1696 3129
rect -1644 3077 -1632 3129
rect -1580 3077 -1380 3129
rect -1328 3077 -1316 3129
rect -1264 3077 -1064 3129
rect -1012 3077 -1000 3129
rect -948 3077 -748 3129
rect -696 3077 -684 3129
rect -632 3077 -432 3129
rect -380 3077 -368 3129
rect -316 3077 -116 3129
rect -64 3077 -52 3129
rect 0 3077 200 3129
rect 252 3077 264 3129
rect 316 3077 516 3129
rect 568 3077 580 3129
rect 632 3077 832 3129
rect 884 3077 896 3129
rect 948 3077 1148 3129
rect 1200 3077 1212 3129
rect 1264 3077 1464 3129
rect 1516 3077 1528 3129
rect 1580 3077 1780 3129
rect 1832 3077 1844 3129
rect 1896 3077 2096 3129
rect 2148 3077 2160 3129
rect 2212 3077 2399 3129
rect -4362 2996 2399 3077
rect -4362 2700 -4140 2996
rect 2453 2900 2550 3196
rect -4081 2819 2550 2900
rect -4081 2767 -4066 2819
rect -4014 2767 -4002 2819
rect -3950 2767 -3750 2819
rect -3698 2767 -3686 2819
rect -3634 2767 -3434 2819
rect -3382 2767 -3370 2819
rect -3318 2767 -3118 2819
rect -3066 2767 -3054 2819
rect -3002 2767 -2802 2819
rect -2750 2767 -2738 2819
rect -2686 2767 -2486 2819
rect -2434 2767 -2422 2819
rect -2370 2767 -2170 2819
rect -2118 2767 -2106 2819
rect -2054 2767 -1854 2819
rect -1802 2767 -1790 2819
rect -1738 2767 -1538 2819
rect -1486 2767 -1474 2819
rect -1422 2767 -1222 2819
rect -1170 2767 -1158 2819
rect -1106 2767 -906 2819
rect -854 2767 -842 2819
rect -790 2767 -590 2819
rect -538 2767 -526 2819
rect -474 2767 -274 2819
rect -222 2767 -210 2819
rect -158 2767 42 2819
rect 94 2767 106 2819
rect 158 2767 358 2819
rect 410 2767 422 2819
rect 474 2767 674 2819
rect 726 2767 738 2819
rect 790 2767 990 2819
rect 1042 2767 1054 2819
rect 1106 2767 1306 2819
rect 1358 2767 1370 2819
rect 1422 2767 1622 2819
rect 1674 2767 1686 2819
rect 1738 2767 1938 2819
rect 1990 2767 2002 2819
rect 2054 2767 2254 2819
rect 2306 2767 2318 2819
rect 2370 2767 2550 2819
rect -4081 2761 2550 2767
rect -4362 2694 2399 2700
rect -4362 2642 -3908 2694
rect -3856 2642 -3844 2694
rect -3792 2642 -3592 2694
rect -3540 2642 -3528 2694
rect -3476 2642 -3276 2694
rect -3224 2642 -3212 2694
rect -3160 2642 -2960 2694
rect -2908 2642 -2896 2694
rect -2844 2642 -2644 2694
rect -2592 2642 -2580 2694
rect -2528 2642 -2328 2694
rect -2276 2642 -2264 2694
rect -2212 2642 -2012 2694
rect -1960 2642 -1948 2694
rect -1896 2642 -1696 2694
rect -1644 2642 -1632 2694
rect -1580 2642 -1380 2694
rect -1328 2642 -1316 2694
rect -1264 2642 -1064 2694
rect -1012 2642 -1000 2694
rect -948 2642 -748 2694
rect -696 2642 -684 2694
rect -632 2642 -432 2694
rect -380 2642 -368 2694
rect -316 2642 -116 2694
rect -64 2642 -52 2694
rect 0 2642 200 2694
rect 252 2642 264 2694
rect 316 2642 516 2694
rect 568 2642 580 2694
rect 632 2642 832 2694
rect 884 2642 896 2694
rect 948 2642 1148 2694
rect 1200 2642 1212 2694
rect 1264 2642 1464 2694
rect 1516 2642 1528 2694
rect 1580 2642 1780 2694
rect 1832 2642 1844 2694
rect 1896 2642 2096 2694
rect 2148 2642 2160 2694
rect 2212 2642 2399 2694
rect -4362 2561 2399 2642
rect -4362 2265 -4140 2561
rect 2453 2465 2550 2761
rect -4081 2384 2550 2465
rect -4081 2332 -4066 2384
rect -4014 2332 -4002 2384
rect -3950 2332 -3750 2384
rect -3698 2332 -3686 2384
rect -3634 2332 -3434 2384
rect -3382 2332 -3370 2384
rect -3318 2332 -3118 2384
rect -3066 2332 -3054 2384
rect -3002 2332 -2802 2384
rect -2750 2332 -2738 2384
rect -2686 2332 -2486 2384
rect -2434 2332 -2422 2384
rect -2370 2332 -2170 2384
rect -2118 2332 -2106 2384
rect -2054 2332 -1854 2384
rect -1802 2332 -1790 2384
rect -1738 2332 -1538 2384
rect -1486 2332 -1474 2384
rect -1422 2332 -1222 2384
rect -1170 2332 -1158 2384
rect -1106 2332 -906 2384
rect -854 2332 -842 2384
rect -790 2332 -590 2384
rect -538 2332 -526 2384
rect -474 2332 -274 2384
rect -222 2332 -210 2384
rect -158 2332 42 2384
rect 94 2332 106 2384
rect 158 2332 358 2384
rect 410 2332 422 2384
rect 474 2332 674 2384
rect 726 2332 738 2384
rect 790 2332 990 2384
rect 1042 2332 1054 2384
rect 1106 2332 1306 2384
rect 1358 2332 1370 2384
rect 1422 2332 1622 2384
rect 1674 2332 1686 2384
rect 1738 2332 1938 2384
rect 1990 2332 2002 2384
rect 2054 2332 2254 2384
rect 2306 2332 2318 2384
rect 2370 2332 2550 2384
rect -4081 2326 2550 2332
rect -4362 2259 2399 2265
rect -4362 2207 -3908 2259
rect -3856 2207 -3844 2259
rect -3792 2207 -3592 2259
rect -3540 2207 -3528 2259
rect -3476 2207 -3276 2259
rect -3224 2207 -3212 2259
rect -3160 2207 -2960 2259
rect -2908 2207 -2896 2259
rect -2844 2207 -2644 2259
rect -2592 2207 -2580 2259
rect -2528 2207 -2328 2259
rect -2276 2207 -2264 2259
rect -2212 2207 -2012 2259
rect -1960 2207 -1948 2259
rect -1896 2207 -1696 2259
rect -1644 2207 -1632 2259
rect -1580 2207 -1380 2259
rect -1328 2207 -1316 2259
rect -1264 2207 -1064 2259
rect -1012 2207 -1000 2259
rect -948 2207 -748 2259
rect -696 2207 -684 2259
rect -632 2207 -432 2259
rect -380 2207 -368 2259
rect -316 2207 -116 2259
rect -64 2207 -52 2259
rect 0 2207 200 2259
rect 252 2207 264 2259
rect 316 2207 516 2259
rect 568 2207 580 2259
rect 632 2207 832 2259
rect 884 2207 896 2259
rect 948 2207 1148 2259
rect 1200 2207 1212 2259
rect 1264 2207 1464 2259
rect 1516 2207 1528 2259
rect 1580 2207 1780 2259
rect 1832 2207 1844 2259
rect 1896 2207 2096 2259
rect 2148 2207 2160 2259
rect 2212 2207 2399 2259
rect -4362 2126 2399 2207
rect -4362 1830 -4140 2126
rect 2453 2030 2550 2326
rect -4081 1949 2550 2030
rect -4081 1897 -4066 1949
rect -4014 1897 -4002 1949
rect -3950 1897 -3750 1949
rect -3698 1897 -3686 1949
rect -3634 1897 -3434 1949
rect -3382 1897 -3370 1949
rect -3318 1897 -3118 1949
rect -3066 1897 -3054 1949
rect -3002 1897 -2802 1949
rect -2750 1897 -2738 1949
rect -2686 1897 -2486 1949
rect -2434 1897 -2422 1949
rect -2370 1897 -2170 1949
rect -2118 1897 -2106 1949
rect -2054 1897 -1854 1949
rect -1802 1897 -1790 1949
rect -1738 1897 -1538 1949
rect -1486 1897 -1474 1949
rect -1422 1897 -1222 1949
rect -1170 1897 -1158 1949
rect -1106 1897 -906 1949
rect -854 1897 -842 1949
rect -790 1897 -590 1949
rect -538 1897 -526 1949
rect -474 1897 -274 1949
rect -222 1897 -210 1949
rect -158 1897 42 1949
rect 94 1897 106 1949
rect 158 1897 358 1949
rect 410 1897 422 1949
rect 474 1897 674 1949
rect 726 1897 738 1949
rect 790 1897 990 1949
rect 1042 1897 1054 1949
rect 1106 1897 1306 1949
rect 1358 1897 1370 1949
rect 1422 1897 1622 1949
rect 1674 1897 1686 1949
rect 1738 1897 1938 1949
rect 1990 1897 2002 1949
rect 2054 1897 2254 1949
rect 2306 1897 2318 1949
rect 2370 1897 2550 1949
rect -4081 1891 2550 1897
rect -4362 1824 2399 1830
rect -4362 1772 -3908 1824
rect -3856 1772 -3844 1824
rect -3792 1772 -3592 1824
rect -3540 1772 -3528 1824
rect -3476 1772 -3276 1824
rect -3224 1772 -3212 1824
rect -3160 1772 -2960 1824
rect -2908 1772 -2896 1824
rect -2844 1772 -2644 1824
rect -2592 1772 -2580 1824
rect -2528 1772 -2328 1824
rect -2276 1772 -2264 1824
rect -2212 1772 -2012 1824
rect -1960 1772 -1948 1824
rect -1896 1772 -1696 1824
rect -1644 1772 -1632 1824
rect -1580 1772 -1380 1824
rect -1328 1772 -1316 1824
rect -1264 1772 -1064 1824
rect -1012 1772 -1000 1824
rect -948 1772 -748 1824
rect -696 1772 -684 1824
rect -632 1772 -432 1824
rect -380 1772 -368 1824
rect -316 1772 -116 1824
rect -64 1772 -52 1824
rect 0 1772 200 1824
rect 252 1772 264 1824
rect 316 1772 516 1824
rect 568 1772 580 1824
rect 632 1772 832 1824
rect 884 1772 896 1824
rect 948 1772 1148 1824
rect 1200 1772 1212 1824
rect 1264 1772 1464 1824
rect 1516 1772 1528 1824
rect 1580 1772 1780 1824
rect 1832 1772 1844 1824
rect 1896 1772 2096 1824
rect 2148 1772 2160 1824
rect 2212 1772 2399 1824
rect -4362 1691 2399 1772
rect -4362 1445 -4140 1691
rect 2453 1508 2550 1891
rect 2666 1508 2683 6104
rect -4362 1402 2363 1445
rect -4362 1401 2147 1402
rect -4362 1400 -3173 1401
rect -4362 1220 -4036 1400
rect -3856 1221 -3173 1400
rect 1295 1222 2147 1401
rect 2327 1222 2363 1402
rect 1295 1221 2363 1222
rect -3856 1220 2363 1221
rect -4362 1177 2363 1220
rect -4362 1176 -4140 1177
rect -4362 932 -4343 1176
rect -4163 932 -4140 1176
rect -4362 911 -4140 932
rect -783 833 821 847
rect -783 832 735 833
rect -4144 779 -3762 789
rect -4144 599 -4098 779
rect -3854 599 -3762 779
rect -783 780 -592 832
rect -540 830 735 832
rect -540 780 -7 830
rect -783 778 -7 780
rect 45 778 415 830
rect 467 781 735 830
rect 787 781 821 833
rect 467 778 821 781
rect -783 769 821 778
rect -783 768 735 769
rect -783 716 -592 768
rect -540 766 735 768
rect -540 716 -7 766
rect -783 714 -7 716
rect 45 714 415 766
rect 467 717 735 766
rect 787 717 821 769
rect 467 714 821 717
rect -783 705 821 714
rect -783 704 735 705
rect -783 652 -592 704
rect -540 702 735 704
rect -540 652 -7 702
rect -783 650 -7 652
rect 45 650 415 702
rect 467 653 735 702
rect 787 653 821 705
rect 467 650 821 653
rect 977 798 1082 1177
rect 977 746 1003 798
rect 1055 746 1082 798
rect 977 734 1082 746
rect 977 682 1003 734
rect 1055 682 1082 734
rect 977 652 1082 682
rect 2453 1002 2683 1508
rect 2453 694 2550 1002
rect 2666 694 2683 1002
rect -783 637 821 650
rect -4144 589 -3762 599
rect -3826 373 -3762 589
rect 2453 633 2683 694
rect 2453 588 2699 633
rect -3705 489 -2097 491
rect -3705 437 -3672 489
rect -3620 437 -3608 489
rect -3556 437 -2507 489
rect -2455 437 -2443 489
rect -2391 437 -2379 489
rect -2327 437 -2315 489
rect -2263 437 -2251 489
rect -2199 437 -2187 489
rect -2135 437 -2097 489
rect -3705 436 -2097 437
rect -1377 487 1975 489
rect -1377 435 -1338 487
rect -1286 435 -1274 487
rect -1222 435 -1210 487
rect -1158 435 -1146 487
rect -1094 435 -1082 487
rect -1030 435 -1018 487
rect -966 435 1755 487
rect 1807 435 1819 487
rect 1871 435 1883 487
rect 1935 435 1975 487
rect -1377 434 1975 435
rect 2453 408 2478 588
rect 2658 408 2699 588
rect -2795 373 -2777 375
rect -3826 323 -2777 373
rect -2725 323 -2713 375
rect -2661 373 -2642 375
rect -1495 373 -1477 375
rect -2661 323 -1477 373
rect -1425 323 -1413 375
rect -1361 373 -1342 375
rect -665 373 -654 375
rect -1361 323 -654 373
rect -602 323 -590 375
rect -538 323 -526 375
rect -474 323 -461 375
rect -3829 213 -3774 235
rect -3228 227 -3210 279
rect -3158 227 -3146 279
rect -3094 277 -3075 279
rect -1927 277 -1909 279
rect -3094 227 -1909 277
rect -1857 227 -1845 279
rect -1793 277 -1774 279
rect -86 277 -75 279
rect -1793 227 -75 277
rect -23 227 -11 279
rect 41 227 53 279
rect 105 277 116 279
rect 2453 277 2699 408
rect 105 227 2699 277
rect -3829 161 -3828 213
rect -3776 174 -3774 213
rect -3776 161 1599 174
rect -3829 149 1599 161
rect -3829 97 -3828 149
rect -3776 132 1599 149
rect -3776 97 -3774 132
rect 1583 122 1599 132
rect 1651 122 1663 174
rect 1715 122 1732 174
rect -3829 76 -3774 97
rect 2453 98 2699 227
rect -4392 1 -4121 44
rect -2293 28 -2264 80
rect -2212 70 -2186 80
rect -987 70 -961 80
rect -2212 28 -961 70
rect -909 70 -883 80
rect 1458 70 1529 78
rect -909 59 1529 70
rect -909 28 1467 59
rect -4392 -307 -4344 1
rect -4164 -307 -4121 1
rect -3221 -67 -2118 -60
rect -3221 -70 -2178 -67
rect -3221 -122 -3214 -70
rect -3162 -122 -2776 -70
rect -2724 -119 -2178 -70
rect -2126 -119 -2118 -67
rect -2724 -122 -2118 -119
rect -3221 -131 -2118 -122
rect -3221 -134 -2178 -131
rect -3221 -186 -3214 -134
rect -3162 -186 -2776 -134
rect -2724 -183 -2178 -134
rect -2126 -183 -2118 -131
rect -2724 -186 -2118 -183
rect -3221 -195 -2118 -186
rect -3221 -198 -2178 -195
rect -3221 -250 -3214 -198
rect -3162 -250 -2776 -198
rect -2724 -247 -2178 -198
rect -2126 -247 -2118 -195
rect -2724 -250 -2118 -247
rect -3221 -256 -2118 -250
rect -1916 -67 -816 -60
rect -1916 -68 -1478 -67
rect -1916 -120 -1907 -68
rect -1855 -119 -1478 -68
rect -1426 -119 -874 -67
rect -822 -119 -816 -67
rect -1855 -120 -816 -119
rect -1916 -131 -816 -120
rect -1916 -132 -1478 -131
rect -1916 -184 -1907 -132
rect -1855 -183 -1478 -132
rect -1426 -183 -874 -131
rect -822 -183 -816 -131
rect -1855 -184 -816 -183
rect -1916 -195 -816 -184
rect -1916 -196 -1478 -195
rect -1916 -248 -1907 -196
rect -1855 -247 -1478 -196
rect -1426 -247 -874 -195
rect -822 -247 -816 -195
rect -1855 -248 -816 -247
rect -1916 -256 -816 -248
rect 239 -112 326 -79
rect 239 -164 257 -112
rect 309 -164 326 -112
rect 239 -176 326 -164
rect 239 -228 257 -176
rect 309 -228 326 -176
rect -4392 -531 -4121 -307
rect -3909 -413 -551 -408
rect -3909 -465 -3861 -413
rect -3809 -465 -3797 -413
rect -3745 -465 -694 -413
rect -642 -465 -630 -413
rect -578 -465 -551 -413
rect -3909 -469 -551 -465
rect 239 -531 326 -228
rect 397 -92 485 28
rect 397 -144 415 -92
rect 467 -144 485 -92
rect 397 -156 485 -144
rect 397 -208 415 -156
rect 467 -208 485 -156
rect 397 -243 485 -208
rect 560 -110 647 -72
rect 560 -162 576 -110
rect 628 -162 647 -110
rect 560 -174 647 -162
rect 560 -226 576 -174
rect 628 -226 647 -174
rect 560 -531 647 -226
rect 717 -92 805 28
rect 717 -144 732 -92
rect 784 -144 805 -92
rect 717 -156 805 -144
rect 717 -208 732 -156
rect 784 -208 805 -156
rect 717 -243 805 -208
rect 879 -109 966 -72
rect 879 -161 894 -109
rect 946 -161 966 -109
rect 879 -173 966 -161
rect 879 -225 894 -173
rect 946 -225 966 -173
rect 879 -531 966 -225
rect 1028 -109 1115 28
rect 1458 7 1467 28
rect 1519 7 1529 59
rect 1458 -5 1529 7
rect 1458 -57 1467 -5
rect 1519 -57 1529 -5
rect 1458 -69 1529 -57
rect 1028 -161 1045 -109
rect 1097 -161 1115 -109
rect 1028 -173 1115 -161
rect 1028 -225 1045 -173
rect 1097 -225 1115 -173
rect 1028 -330 1115 -225
rect 1312 -107 1399 -73
rect 1312 -159 1327 -107
rect 1379 -159 1399 -107
rect 1312 -171 1399 -159
rect 1312 -223 1327 -171
rect 1379 -223 1399 -171
rect 1312 -531 1399 -223
rect 1458 -121 1467 -69
rect 1519 -121 1529 -69
rect 1458 -133 1529 -121
rect 1458 -185 1467 -133
rect 1519 -185 1529 -133
rect 1458 -197 1529 -185
rect 1458 -249 1467 -197
rect 1519 -249 1529 -197
rect 1458 -261 1529 -249
rect 1458 -313 1467 -261
rect 1519 -313 1529 -261
rect 1458 -337 1529 -313
rect 2453 -82 2478 98
rect 2658 -82 2699 98
rect -4392 -574 2271 -531
rect -4392 -626 -3657 -574
rect -3605 -626 -3593 -574
rect -3541 -626 -3529 -574
rect -3477 -626 -3465 -574
rect -3413 -626 -3401 -574
rect -3349 -626 -3337 -574
rect -3285 -626 -3273 -574
rect -3221 -626 -3209 -574
rect -3157 -626 -3145 -574
rect -3093 -626 -3081 -574
rect -3029 -626 -3017 -574
rect -2965 -626 -2953 -574
rect -2901 -626 -2889 -574
rect -2837 -626 -2825 -574
rect -2773 -626 -2761 -574
rect -2709 -626 -2697 -574
rect -2645 -626 -2633 -574
rect -2581 -626 -2569 -574
rect -2517 -626 -2505 -574
rect -2453 -626 -2441 -574
rect -2389 -626 -2377 -574
rect -2325 -626 -2313 -574
rect -2261 -626 -2249 -574
rect -2197 -626 -2185 -574
rect -2133 -626 -2121 -574
rect -2069 -626 -2057 -574
rect -2005 -626 -1993 -574
rect -1941 -626 -1929 -574
rect -1877 -626 -1865 -574
rect -1813 -626 -1801 -574
rect -1749 -626 -1737 -574
rect -1685 -626 -1673 -574
rect -1621 -626 -1609 -574
rect -1557 -626 -1545 -574
rect -1493 -626 -1481 -574
rect -1429 -626 -1417 -574
rect -1365 -626 -1353 -574
rect -1301 -626 -1289 -574
rect -1237 -626 -1225 -574
rect -1173 -626 -1161 -574
rect -1109 -626 -1097 -574
rect -1045 -626 -1033 -574
rect -981 -626 -969 -574
rect -917 -626 -905 -574
rect -853 -626 -841 -574
rect -789 -626 -777 -574
rect -725 -626 -713 -574
rect -661 -626 -649 -574
rect -597 -626 -585 -574
rect -533 -626 -521 -574
rect -469 -626 -457 -574
rect -405 -626 -393 -574
rect -341 -626 -329 -574
rect -277 -626 -265 -574
rect -213 -626 -201 -574
rect -149 -626 -137 -574
rect -85 -626 -73 -574
rect -21 -626 -9 -574
rect 43 -626 55 -574
rect 107 -626 119 -574
rect 171 -626 183 -574
rect 235 -626 247 -574
rect 299 -626 311 -574
rect 363 -626 375 -574
rect 427 -626 439 -574
rect 491 -626 503 -574
rect 555 -626 567 -574
rect 619 -626 631 -574
rect 683 -626 695 -574
rect 747 -626 759 -574
rect 811 -626 823 -574
rect 875 -626 887 -574
rect 939 -626 951 -574
rect 1003 -626 1015 -574
rect 1067 -626 1079 -574
rect 1131 -626 1143 -574
rect 1195 -626 1207 -574
rect 1259 -626 1271 -574
rect 1323 -626 1335 -574
rect 1387 -626 1399 -574
rect 1451 -626 1463 -574
rect 1515 -626 1527 -574
rect 1579 -626 1591 -574
rect 1643 -626 1655 -574
rect 1707 -626 1719 -574
rect 1771 -626 1783 -574
rect 1835 -626 1847 -574
rect 1899 -626 1911 -574
rect 1963 -626 1975 -574
rect 2027 -626 2039 -574
rect 2091 -626 2103 -574
rect 2155 -626 2167 -574
rect 2219 -626 2271 -574
rect -4392 -685 2271 -626
rect -4392 -1003 -4121 -685
rect 2453 -803 2699 -82
rect -4092 -884 2699 -803
rect -4092 -936 -4066 -884
rect -4014 -936 -4002 -884
rect -3950 -936 -3750 -884
rect -3698 -936 -3686 -884
rect -3634 -936 -3434 -884
rect -3382 -936 -3370 -884
rect -3318 -936 -3118 -884
rect -3066 -936 -3054 -884
rect -3002 -936 -2802 -884
rect -2750 -936 -2738 -884
rect -2686 -936 -2486 -884
rect -2434 -936 -2422 -884
rect -2370 -936 -2170 -884
rect -2118 -936 -2106 -884
rect -2054 -936 -1854 -884
rect -1802 -936 -1790 -884
rect -1738 -936 -1538 -884
rect -1486 -936 -1474 -884
rect -1422 -936 -1222 -884
rect -1170 -936 -1158 -884
rect -1106 -936 -906 -884
rect -854 -936 -842 -884
rect -790 -936 -590 -884
rect -538 -936 -526 -884
rect -474 -936 -274 -884
rect -222 -936 -210 -884
rect -158 -936 42 -884
rect 94 -936 106 -884
rect 158 -936 358 -884
rect 410 -936 422 -884
rect 474 -936 674 -884
rect 726 -936 738 -884
rect 790 -936 990 -884
rect 1042 -936 1054 -884
rect 1106 -936 1306 -884
rect 1358 -936 1370 -884
rect 1422 -936 1622 -884
rect 1674 -936 1686 -884
rect 1738 -936 1938 -884
rect 1990 -936 2002 -884
rect 2054 -936 2254 -884
rect 2306 -936 2318 -884
rect 2370 -936 2699 -884
rect -4092 -942 2699 -936
rect -4393 -1009 2383 -1003
rect -4393 -1061 -3908 -1009
rect -3856 -1061 -3844 -1009
rect -3792 -1061 -3592 -1009
rect -3540 -1061 -3528 -1009
rect -3476 -1061 -3276 -1009
rect -3224 -1061 -3212 -1009
rect -3160 -1061 -2960 -1009
rect -2908 -1061 -2896 -1009
rect -2844 -1061 -2644 -1009
rect -2592 -1061 -2580 -1009
rect -2528 -1061 -2328 -1009
rect -2276 -1061 -2264 -1009
rect -2212 -1061 -2012 -1009
rect -1960 -1061 -1948 -1009
rect -1896 -1061 -1696 -1009
rect -1644 -1061 -1632 -1009
rect -1580 -1061 -1380 -1009
rect -1328 -1061 -1316 -1009
rect -1264 -1061 -1064 -1009
rect -1012 -1061 -1000 -1009
rect -948 -1061 -748 -1009
rect -696 -1061 -684 -1009
rect -632 -1061 -432 -1009
rect -380 -1061 -368 -1009
rect -316 -1061 -116 -1009
rect -64 -1061 -52 -1009
rect 0 -1061 200 -1009
rect 252 -1061 264 -1009
rect 316 -1061 516 -1009
rect 568 -1061 580 -1009
rect 632 -1061 832 -1009
rect 884 -1061 896 -1009
rect 948 -1061 1148 -1009
rect 1200 -1061 1212 -1009
rect 1264 -1061 1464 -1009
rect 1516 -1061 1528 -1009
rect 1580 -1061 1780 -1009
rect 1832 -1061 1844 -1009
rect 1896 -1061 2096 -1009
rect 2148 -1061 2160 -1009
rect 2212 -1061 2383 -1009
rect -4393 -1142 2383 -1061
rect -4392 -1421 -4121 -1142
rect 2437 -1221 2699 -942
rect -4081 -1302 2699 -1221
rect -4081 -1354 -4066 -1302
rect -4014 -1354 -4002 -1302
rect -3950 -1354 -3750 -1302
rect -3698 -1354 -3686 -1302
rect -3634 -1354 -3434 -1302
rect -3382 -1354 -3370 -1302
rect -3318 -1354 -3118 -1302
rect -3066 -1354 -3054 -1302
rect -3002 -1354 -2802 -1302
rect -2750 -1354 -2738 -1302
rect -2686 -1354 -2486 -1302
rect -2434 -1354 -2422 -1302
rect -2370 -1354 -2170 -1302
rect -2118 -1354 -2106 -1302
rect -2054 -1354 -1854 -1302
rect -1802 -1354 -1790 -1302
rect -1738 -1354 -1538 -1302
rect -1486 -1354 -1474 -1302
rect -1422 -1354 -1222 -1302
rect -1170 -1354 -1158 -1302
rect -1106 -1354 -906 -1302
rect -854 -1354 -842 -1302
rect -790 -1354 -590 -1302
rect -538 -1354 -526 -1302
rect -474 -1354 -274 -1302
rect -222 -1354 -210 -1302
rect -158 -1354 42 -1302
rect 94 -1354 106 -1302
rect 158 -1354 358 -1302
rect 410 -1354 422 -1302
rect 474 -1354 674 -1302
rect 726 -1354 738 -1302
rect 790 -1354 990 -1302
rect 1042 -1354 1054 -1302
rect 1106 -1354 1306 -1302
rect 1358 -1354 1370 -1302
rect 1422 -1354 1622 -1302
rect 1674 -1354 1686 -1302
rect 1738 -1354 1938 -1302
rect 1990 -1354 2002 -1302
rect 2054 -1354 2254 -1302
rect 2306 -1354 2318 -1302
rect 2370 -1354 2699 -1302
rect -4081 -1360 2699 -1354
rect -4392 -1427 2383 -1421
rect -4392 -1479 -3908 -1427
rect -3856 -1479 -3844 -1427
rect -3792 -1479 -3592 -1427
rect -3540 -1479 -3528 -1427
rect -3476 -1479 -3276 -1427
rect -3224 -1479 -3212 -1427
rect -3160 -1479 -2960 -1427
rect -2908 -1479 -2896 -1427
rect -2844 -1479 -2644 -1427
rect -2592 -1479 -2580 -1427
rect -2528 -1479 -2328 -1427
rect -2276 -1479 -2264 -1427
rect -2212 -1479 -2012 -1427
rect -1960 -1479 -1948 -1427
rect -1896 -1479 -1696 -1427
rect -1644 -1479 -1632 -1427
rect -1580 -1479 -1380 -1427
rect -1328 -1479 -1316 -1427
rect -1264 -1479 -1064 -1427
rect -1012 -1479 -1000 -1427
rect -948 -1479 -748 -1427
rect -696 -1479 -684 -1427
rect -632 -1479 -432 -1427
rect -380 -1479 -368 -1427
rect -316 -1479 -116 -1427
rect -64 -1479 -52 -1427
rect 0 -1479 200 -1427
rect 252 -1479 264 -1427
rect 316 -1479 516 -1427
rect 568 -1479 580 -1427
rect 632 -1479 832 -1427
rect 884 -1479 896 -1427
rect 948 -1479 1148 -1427
rect 1200 -1479 1212 -1427
rect 1264 -1479 1464 -1427
rect 1516 -1479 1528 -1427
rect 1580 -1479 1780 -1427
rect 1832 -1479 1844 -1427
rect 1896 -1479 2096 -1427
rect 2148 -1479 2160 -1427
rect 2212 -1479 2383 -1427
rect -4392 -1560 2383 -1479
rect -4392 -1839 -4121 -1560
rect 2437 -1639 2699 -1360
rect -4081 -1720 2699 -1639
rect -4081 -1772 -4066 -1720
rect -4014 -1772 -4002 -1720
rect -3950 -1772 -3750 -1720
rect -3698 -1772 -3686 -1720
rect -3634 -1772 -3434 -1720
rect -3382 -1772 -3370 -1720
rect -3318 -1772 -3118 -1720
rect -3066 -1772 -3054 -1720
rect -3002 -1772 -2802 -1720
rect -2750 -1772 -2738 -1720
rect -2686 -1772 -2486 -1720
rect -2434 -1772 -2422 -1720
rect -2370 -1772 -2170 -1720
rect -2118 -1772 -2106 -1720
rect -2054 -1772 -1854 -1720
rect -1802 -1772 -1790 -1720
rect -1738 -1772 -1538 -1720
rect -1486 -1772 -1474 -1720
rect -1422 -1772 -1222 -1720
rect -1170 -1772 -1158 -1720
rect -1106 -1772 -906 -1720
rect -854 -1772 -842 -1720
rect -790 -1772 -590 -1720
rect -538 -1772 -526 -1720
rect -474 -1772 -274 -1720
rect -222 -1772 -210 -1720
rect -158 -1772 42 -1720
rect 94 -1772 106 -1720
rect 158 -1772 358 -1720
rect 410 -1772 422 -1720
rect 474 -1772 674 -1720
rect 726 -1772 738 -1720
rect 790 -1772 990 -1720
rect 1042 -1772 1054 -1720
rect 1106 -1772 1306 -1720
rect 1358 -1772 1370 -1720
rect 1422 -1772 1622 -1720
rect 1674 -1772 1686 -1720
rect 1738 -1772 1938 -1720
rect 1990 -1772 2002 -1720
rect 2054 -1772 2254 -1720
rect 2306 -1772 2318 -1720
rect 2370 -1772 2699 -1720
rect -4081 -1778 2699 -1772
rect -4392 -1845 2383 -1839
rect -4392 -1897 -3908 -1845
rect -3856 -1897 -3844 -1845
rect -3792 -1897 -3592 -1845
rect -3540 -1897 -3528 -1845
rect -3476 -1897 -3276 -1845
rect -3224 -1897 -3212 -1845
rect -3160 -1897 -2960 -1845
rect -2908 -1897 -2896 -1845
rect -2844 -1897 -2644 -1845
rect -2592 -1897 -2580 -1845
rect -2528 -1897 -2328 -1845
rect -2276 -1897 -2264 -1845
rect -2212 -1897 -2012 -1845
rect -1960 -1897 -1948 -1845
rect -1896 -1897 -1696 -1845
rect -1644 -1897 -1632 -1845
rect -1580 -1897 -1380 -1845
rect -1328 -1897 -1316 -1845
rect -1264 -1897 -1064 -1845
rect -1012 -1897 -1000 -1845
rect -948 -1897 -748 -1845
rect -696 -1897 -684 -1845
rect -632 -1897 -432 -1845
rect -380 -1897 -368 -1845
rect -316 -1897 -116 -1845
rect -64 -1897 -52 -1845
rect 0 -1897 200 -1845
rect 252 -1897 264 -1845
rect 316 -1897 516 -1845
rect 568 -1897 580 -1845
rect 632 -1897 832 -1845
rect 884 -1897 896 -1845
rect 948 -1897 1148 -1845
rect 1200 -1897 1212 -1845
rect 1264 -1897 1464 -1845
rect 1516 -1897 1528 -1845
rect 1580 -1897 1780 -1845
rect 1832 -1897 1844 -1845
rect 1896 -1897 2096 -1845
rect 2148 -1897 2160 -1845
rect 2212 -1897 2383 -1845
rect -4392 -1978 2383 -1897
rect -4392 -2131 -4121 -1978
rect -4392 -2439 -4380 -2131
rect -4136 -2439 -4121 -2131
rect -4392 -2472 -4121 -2439
rect 1573 -3234 2705 -3220
rect 1573 -3286 2638 -3234
rect 2690 -3286 2705 -3234
rect 1573 -3296 2705 -3286
rect 1573 -3412 1631 -3296
rect 2195 -3298 2705 -3296
rect 2195 -3350 2638 -3298
rect 2690 -3350 2705 -3298
rect 2195 -3362 2705 -3350
rect 2195 -3412 2638 -3362
rect 1573 -3414 2638 -3412
rect 2690 -3414 2705 -3362
rect 1573 -3426 2705 -3414
rect 1573 -3478 2638 -3426
rect 2690 -3478 2705 -3426
rect 1573 -3491 2705 -3478
use sky130_fd_pr__nfet_g5v0d10v5_EJGQJV  M13
timestamp 1694031861
transform 1 0 1710 0 1 -157
box -268 -348 268 348
use sky130_fd_pr__nfet_g5v0d10v5_EJGQJV  M24
timestamp 1694031861
transform 1 0 1275 0 1 -157
box -268 -348 268 348
use sky130_fd_pr__diode_pw2nd_05v5_L93GHW  sky130_fd_pr__diode_pw2nd_05v5_L93GHW_0
timestamp 1694031861
transform 1 0 -3804 0 1 -100
box -188 -188 188 188
use sky130_fd_pr__diode_pw2nd_05v5_L93GHW  sky130_fd_pr__diode_pw2nd_05v5_L93GHW_1
timestamp 1694031861
transform 1 0 -3804 0 1 500
box -188 -188 188 188
use sky130_fd_pr__nfet_03v3_nvt_EJGQJV  sky130_fd_pr__nfet_03v3_nvt_EJGQJV_0
timestamp 1694031861
transform -1 0 -2671 0 1 -157
box -268 -348 268 348
use sky130_fd_pr__pfet_g5v0d10v5_AQ2AJT  sky130_fd_pr__pfet_g5v0d10v5_AQ2AJT_0
timestamp 1694031861
transform 1 0 -849 0 1 2735
box -3389 -1269 3389 1269
use sky130_fd_pr__pfet_g5v0d10v5_AQ2AJT  sky130_fd_pr__pfet_g5v0d10v5_AQ2AJT_1
timestamp 1694031861
transform 1 0 -849 0 1 5083
box -3389 -1269 3389 1269
use sky130_fd_pr__res_xhigh_po_0p35_D7NTZ8  sky130_fd_pr__res_xhigh_po_0p35_D7NTZ8_0
timestamp 1694031861
transform 0 1 -890 -1 0 -2878
box -668 -3088 668 3088
use sky130_fd_pr__nfet_g5v0d10v5_EJGQJV  XM1
timestamp 1694031861
transform -1 0 -1803 0 1 -157
box -268 -348 268 348
use sky130_fd_pr__nfet_g5v0d10v5_EJGQJV  XM2
timestamp 1694031861
transform -1 0 -1369 0 1 -157
box -268 -348 268 348
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  XM3
timestamp 1694031861
transform 1 0 -2319 0 1 704
box -387 -362 387 362
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  XM4
timestamp 1694031861
transform -1 0 -1151 0 1 704
box -387 -362 387 362
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  XM5
timestamp 1694031861
transform -1 0 -1735 0 1 704
box -387 -362 387 362
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  XM6
timestamp 1694031861
transform 1 0 -2903 0 1 704
box -387 -362 387 362
use sky130_fd_pr__nfet_g5v0d10v5_EJGQJV  XM7
timestamp 1694031861
transform -1 0 -2237 0 1 -157
box -268 -348 268 348
use sky130_fd_pr__nfet_03v3_nvt_EJGQJV  XM8
timestamp 1694031861
transform -1 0 -3105 0 1 -157
box -268 -348 268 348
use sky130_fd_pr__nfet_g5v0d10v5_EJGQJV  XM9
timestamp 1694031861
transform -1 0 -935 0 1 -157
box -268 -348 268 348
use sky130_fd_pr__nfet_g5v0d10v5_H7BQ24  XM10
timestamp 1694031861
transform 1 0 603 0 1 -158
box -505 -348 505 348
use sky130_fd_pr__nfet_g5v0d10v5_UC3VEF  XM22
timestamp 1694031861
transform 1 0 -865 0 1 -1392
box -3349 -766 3349 766
use sky130_fd_pr__pfet_g5v0d10v5_U6NWY6  XM25
timestamp 1694031861
transform 1 0 1106 0 1 704
box -308 -362 308 362
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  XM26
timestamp 1694031861
transform 1 0 601 0 1 704
box -387 -362 387 362
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  XM27
timestamp 1694031861
transform 1 0 17 0 1 704
box -387 -362 387 362
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  XM28
timestamp 1694031861
transform 1 0 -567 0 1 704
box -387 -362 387 362
use sky130_fd_pr__nfet_g5v0d10v5_EJGQJV  XM29
timestamp 1694031861
transform -1 0 -501 0 1 -157
box -268 -348 268 348
use sky130_fd_pr__nfet_g5v0d10v5_EJGQJV  XM30
timestamp 1694031861
transform -1 0 -67 0 1 -157
box -268 -348 268 348
<< labels >>
flabel metal2 s -241 738 -241 738 0 FreeSans 256 0 0 0 vcomp
flabel metal2 s -3529 -437 -3529 -437 0 FreeSans 256 0 0 0 ndrv
flabel metal2 s 1374 46 1374 46 0 FreeSans 256 0 0 0 nbias
flabel metal1 s 980 577 980 577 0 FreeSans 256 0 0 0 pbias
flabel metal2 s -3326 462 -3326 462 0 FreeSans 256 0 0 0 pdrv2
flabel metal2 s 1468 463 1468 463 0 FreeSans 256 0 0 0 pdrv1
flabel metal2 s -2456 -160 -2456 -160 0 FreeSans 256 0 0 0 vcomn2
flabel metal2 s -1322 -168 -1322 -168 0 FreeSans 256 0 0 0 vcomn1
flabel metal1 s -4342 1201 -4142 1401 0 FreeSans 205 0 0 0 vdd
port 1 nsew
flabel metal1 s -4361 589 -4161 789 0 FreeSans 205 0 0 0 in
port 2 nsew
flabel metal1 s 2467 163 2667 363 0 FreeSans 205 0 0 0 out
port 3 nsew
flabel metal1 s -4355 -529 -4155 -329 0 FreeSans 205 0 0 0 vss
port 4 nsew
flabel metal1 s -4361 244 -4161 444 0 FreeSans 256 0 0 0 ena
port 5 nsew
<< end >>
