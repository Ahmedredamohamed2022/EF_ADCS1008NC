magic
tech sky130A
magscale 1 2
timestamp 1699205827
<< checkpaint >>
rect -2810 -93421 68824 14266
<< metal1 >>
rect -422 96 112 122
rect -422 64 -409 96
rect -426 -20 -409 64
rect 91 64 112 96
rect 91 -20 1080 64
rect -426 -40 1080 -20
rect 596 -2746 1002 -2721
rect 596 -2990 613 -2746
rect 985 -2990 1002 -2746
rect 596 -3015 1002 -2990
rect -1199 -3549 158 -3544
rect -1199 -3571 164 -3549
rect -1199 -3687 -1173 -3571
rect -609 -3687 164 -3571
rect -1199 -3746 164 -3687
rect -36 -3749 164 -3746
rect 210 -6227 492 -6203
rect 210 -6471 229 -6227
rect 473 -6471 492 -6227
rect 210 -6495 492 -6471
rect 1806 -6687 2106 -6641
rect 1806 -7315 1838 -6687
rect 2082 -7315 2106 -6687
rect 1806 -7375 2106 -7315
rect -420 -7514 164 -7469
rect -420 -7630 -385 -7514
rect 115 -7630 164 -7514
rect -420 -7667 164 -7630
rect -398 -7669 164 -7667
rect 33370 -7790 33860 -7782
rect -42 -7814 164 -7805
rect -404 -7848 240 -7814
rect -404 -7964 -366 -7848
rect 198 -7964 240 -7848
rect 32094 -7828 33860 -7790
rect 19858 -7882 20052 -7878
rect -404 -7998 240 -7964
rect 19296 -7921 20052 -7882
rect -42 -8015 164 -7998
rect 19296 -8037 19899 -7921
rect 20015 -8037 20052 -7921
rect 19296 -8080 20052 -8037
rect 19300 -8081 19432 -8080
rect 32094 -8136 33429 -7828
rect 33801 -8136 33860 -7828
rect 32094 -8198 33860 -8136
<< via1 >>
rect -409 -20 91 96
rect 613 -2990 985 -2746
rect -1173 -3687 -609 -3571
rect 229 -6471 473 -6227
rect 1838 -7315 2082 -6687
rect -385 -7630 115 -7514
rect -366 -7964 198 -7848
rect 19899 -8037 20015 -7921
rect 33429 -8136 33801 -7828
<< metal2 >>
rect 3218 12706 3310 13002
rect 6616 12702 6708 12998
rect 10014 12702 10106 12998
rect 13318 12700 13410 12996
rect 16628 12706 16720 13002
rect 20004 12702 20100 13004
rect 23308 12698 23404 13000
rect 26752 12698 26843 12996
rect 26672 8732 26930 8788
rect 26672 8514 26689 8732
rect 26660 8276 26689 8514
rect 26905 8276 26930 8732
rect 26660 8214 26930 8276
rect 26660 8016 26922 8214
rect -422 106 112 122
rect -422 96 -387 106
rect 69 96 112 106
rect -422 -20 -409 96
rect 91 -20 112 96
rect -422 -30 -387 -20
rect 69 -30 112 -20
rect -422 -40 112 -30
rect 576 -114 912 -104
rect 576 -170 595 -114
rect 651 -170 675 -114
rect 731 -170 755 -114
rect 811 -170 835 -114
rect 891 -170 912 -114
rect 200 -293 510 -273
rect 200 -349 245 -293
rect 301 -349 325 -293
rect 381 -349 405 -293
rect 461 -349 510 -293
rect 200 -2701 510 -349
rect 198 -3031 510 -2701
rect -1208 -3561 -578 -3532
rect -1208 -3571 -1159 -3561
rect -623 -3571 -578 -3561
rect -1208 -3687 -1173 -3571
rect -609 -3687 -578 -3571
rect -1208 -3697 -1159 -3687
rect -623 -3697 -578 -3687
rect -1208 -3734 -578 -3697
rect 200 -6227 510 -3031
rect 576 -2385 912 -170
rect 26700 -288 26922 8016
rect 26700 -344 26740 -288
rect 26796 -344 26820 -288
rect 26876 -344 26922 -288
rect 26700 -365 26922 -344
rect 1802 -480 2102 -436
rect 1802 -776 1843 -480
rect 2059 -776 2102 -480
rect 576 -2699 1030 -2385
rect 576 -2746 1036 -2699
rect 576 -2990 613 -2746
rect 985 -2990 1036 -2746
rect 576 -3049 1036 -2990
rect 200 -6471 229 -6227
rect 473 -6471 510 -6227
rect 200 -6500 510 -6471
rect 1802 -6641 2102 -776
rect 1802 -6687 2106 -6641
rect 1802 -7315 1838 -6687
rect 2082 -7315 2106 -6687
rect 1802 -7349 2106 -7315
rect 1806 -7375 2106 -7349
rect -420 -7504 164 -7469
rect -420 -7514 -363 -7504
rect 93 -7514 164 -7504
rect -420 -7630 -385 -7514
rect 115 -7630 164 -7514
rect -420 -7640 -363 -7630
rect 93 -7640 164 -7630
rect -420 -7667 164 -7640
rect -404 -7838 240 -7814
rect -404 -7848 -352 -7838
rect 184 -7848 240 -7838
rect -404 -7964 -366 -7848
rect 198 -7964 240 -7848
rect 33370 -7828 33860 -7782
rect 33370 -7834 33429 -7828
rect 33801 -7834 33860 -7828
rect -404 -7974 -352 -7964
rect 184 -7974 240 -7964
rect -404 -7998 240 -7974
rect 19858 -7911 20052 -7878
rect 19858 -8047 19889 -7911
rect 20025 -8047 20052 -7911
rect 19858 -8078 20052 -8047
rect 33370 -8130 33427 -7834
rect 33803 -8130 33860 -7834
rect 33370 -8136 33429 -8130
rect 33801 -8136 33860 -8130
rect 33370 -8190 33860 -8136
rect 32420 -10343 32596 -10214
rect 32420 -10479 32437 -10343
rect 32573 -10479 32596 -10343
rect 32420 -10510 32596 -10479
rect 17992 -13291 18604 -13206
rect 17992 -13747 18095 -13291
rect 18471 -13747 18604 -13291
rect 17992 -13816 18604 -13747
rect 18136 -14740 18400 -13816
rect 22384 -14248 23000 -14180
rect 22384 -14704 22449 -14248
rect 22905 -14704 23000 -14248
rect 30990 -14534 31542 -14532
rect 18164 -15068 18386 -14740
rect 22384 -14774 23000 -14704
rect 30988 -14623 31552 -14534
rect 22560 -15060 22776 -14774
rect 30988 -14999 31042 -14623
rect 31498 -14999 31552 -14623
rect 30988 -15072 31552 -14999
rect 30990 -15090 31542 -15072
rect 31126 -15190 31348 -15090
<< via2 >>
rect 26689 8276 26905 8732
rect -387 96 69 106
rect -387 -20 69 96
rect -387 -30 69 -20
rect 595 -170 651 -114
rect 675 -170 731 -114
rect 755 -170 811 -114
rect 835 -170 891 -114
rect 245 -349 301 -293
rect 325 -349 381 -293
rect 405 -349 461 -293
rect -1159 -3571 -623 -3561
rect -1159 -3687 -623 -3571
rect -1159 -3697 -623 -3687
rect 26740 -344 26796 -288
rect 26820 -344 26876 -288
rect 1843 -776 2059 -480
rect -363 -7514 93 -7504
rect -363 -7630 93 -7514
rect -363 -7640 93 -7630
rect -352 -7848 184 -7838
rect -352 -7964 184 -7848
rect -352 -7974 184 -7964
rect 19889 -7921 20025 -7911
rect 19889 -8037 19899 -7921
rect 19899 -8037 20015 -7921
rect 20015 -8037 20025 -7921
rect 19889 -8047 20025 -8037
rect 33427 -8130 33429 -7834
rect 33429 -8130 33801 -7834
rect 33801 -8130 33803 -7834
rect 32437 -10479 32573 -10343
rect 18095 -13747 18471 -13291
rect 22449 -14704 22905 -14248
rect 31042 -14999 31498 -14623
<< metal3 >>
rect 26672 8736 26930 8788
rect 26672 8272 26685 8736
rect 26909 8272 26930 8736
rect 26672 8214 26930 8272
rect 33702 6816 34010 6876
rect 33700 6678 34008 6738
rect 33704 6544 34012 6604
rect 20094 4278 20302 4318
rect 20094 4214 20125 4278
rect 20189 4214 20205 4278
rect 20269 4214 20302 4278
rect 20094 4166 20302 4214
rect -422 106 112 122
rect -422 70 -387 106
rect 69 70 112 106
rect -422 6 -391 70
rect 73 6 112 70
rect -422 -30 -387 6
rect 69 -30 112 6
rect -422 -40 112 -30
rect 0 -114 35086 -102
rect 0 -170 595 -114
rect 651 -170 675 -114
rect 731 -170 755 -114
rect 811 -170 835 -114
rect 891 -116 35086 -114
rect 891 -170 23448 -116
rect 0 -180 23448 -170
rect 23512 -180 23528 -116
rect 23592 -180 23608 -116
rect 23672 -180 23688 -116
rect 23752 -118 35086 -116
rect 23752 -180 32850 -118
rect 0 -182 32850 -180
rect 32914 -182 32930 -118
rect 32994 -182 33010 -118
rect 33074 -182 33090 -118
rect 33154 -182 35086 -118
rect 0 -196 35086 -182
rect -4 -280 35086 -272
rect -6 -285 35086 -280
rect -6 -288 33384 -285
rect -6 -293 26740 -288
rect -6 -349 245 -293
rect 301 -349 325 -293
rect 381 -349 405 -293
rect 461 -344 26740 -293
rect 26796 -344 26820 -288
rect 26876 -344 33384 -288
rect 461 -349 33384 -344
rect 33448 -349 33464 -285
rect 33528 -349 33544 -285
rect 33608 -349 33624 -285
rect 33688 -349 33704 -285
rect 33768 -349 33784 -285
rect 33848 -349 35086 -285
rect -6 -366 35086 -349
rect -6 -370 292 -366
rect -6 -436 1144 -434
rect -10 -464 35086 -436
rect -10 -480 34037 -464
rect -10 -776 1843 -480
rect 2059 -481 34037 -480
rect 2059 -625 20123 -481
rect 20267 -625 34037 -481
rect 2059 -768 34037 -625
rect 34421 -768 35086 -464
rect 2059 -776 35086 -768
rect -10 -836 35086 -776
rect 0 -958 35086 -918
rect 0 -1228 1059 -958
rect 14 -1262 1059 -1228
rect 1363 -966 35086 -958
rect 1363 -1262 31466 -966
rect 14 -1270 31466 -1262
rect 31610 -973 35086 -966
rect 31610 -1270 34635 -973
rect 14 -1277 34635 -1270
rect 35019 -1277 35086 -973
rect 14 -1318 35086 -1277
rect -1208 -3561 -578 -3544
rect -1208 -3697 -1159 -3561
rect -623 -3697 -578 -3561
rect -1208 -3746 -578 -3697
rect 32400 -7252 33212 -7196
rect -420 -7500 164 -7469
rect -420 -7644 -367 -7500
rect 97 -7644 164 -7500
rect -420 -7667 164 -7644
rect 32400 -7636 32854 -7252
rect 33158 -7636 33212 -7252
rect 32400 -7700 33212 -7636
rect -1208 -7812 -650 -7806
rect -1210 -7814 236 -7812
rect -1210 -7834 240 -7814
rect -1210 -7978 -356 -7834
rect 188 -7978 240 -7834
rect 33370 -7830 33860 -7782
rect -1210 -7992 240 -7978
rect -404 -7998 240 -7992
rect 19858 -7911 20050 -7862
rect 19858 -8047 19889 -7911
rect 20025 -8047 20050 -7911
rect 19858 -9574 20050 -8047
rect 33370 -8134 33423 -7830
rect 33807 -8134 33860 -7830
rect 33370 -8190 33860 -8134
rect 33588 -8296 34002 -8292
rect 31794 -8488 34002 -8296
rect 33588 -8490 34002 -8488
rect 17992 -13291 18604 -13206
rect 17992 -13747 18095 -13291
rect 18471 -13408 18604 -13291
rect 19860 -13408 20052 -9675
rect 32420 -10243 32596 -10214
rect 32420 -10467 32433 -10243
rect 32577 -10467 32596 -10243
rect 32420 -10479 32437 -10467
rect 32573 -10479 32596 -10467
rect 32420 -10510 32596 -10479
rect 18471 -13600 20052 -13408
rect 18471 -13747 18604 -13600
rect 17992 -13816 18604 -13747
rect 22384 -14192 23000 -14180
rect -408 -14196 32280 -14192
rect -408 -14225 32630 -14196
rect -408 -14369 -356 -14225
rect -52 -14248 32630 -14225
rect -52 -14369 22449 -14248
rect -408 -14388 22449 -14369
rect -404 -14392 22449 -14388
rect 22384 -14704 22449 -14392
rect 22905 -14267 32630 -14248
rect 22905 -14331 32238 -14267
rect 32302 -14331 32318 -14267
rect 32382 -14331 32398 -14267
rect 32462 -14331 32478 -14267
rect 32542 -14331 32558 -14267
rect 32622 -14331 32630 -14267
rect 22905 -14392 32630 -14331
rect 22905 -14704 23000 -14392
rect 32200 -14406 32630 -14392
rect 30990 -14534 31542 -14532
rect 22384 -14774 23000 -14704
rect 30988 -14623 31552 -14534
rect -406 -14894 414 -14884
rect 30988 -14894 31042 -14623
rect -406 -14999 31042 -14894
rect 31498 -14999 31552 -14623
rect -406 -15072 31552 -14999
rect -406 -15086 31542 -15072
rect 30990 -15090 31542 -15086
rect 32838 -15296 33164 -15276
rect 32838 -15760 32849 -15296
rect 33153 -15760 33164 -15296
rect 32838 -15780 33164 -15760
rect 33388 -16079 33820 -16078
rect 33388 -16543 33412 -16079
rect 33796 -16543 33820 -16079
rect 33388 -16544 33820 -16543
rect 34048 -16901 34454 -16896
rect 34048 -17365 34059 -16901
rect 34443 -17365 34454 -16901
rect 34048 -17370 34454 -17365
rect 34616 -17704 35036 -17676
rect 34616 -18168 34634 -17704
rect 35018 -18168 35036 -17704
rect 34616 -18196 35036 -18168
rect -6 -26596 1146 -26420
rect -2 -33322 1150 -33146
rect -10 -40038 1142 -39862
rect 2 -46732 1154 -46556
rect 6 -53502 1158 -53326
rect -6 -54414 1146 -54238
rect -16 -54880 1136 -54704
rect -6 -60488 1146 -60312
rect 2 -67194 1154 -67018
rect -2 -73914 1150 -73738
rect -10 -80616 1142 -80440
rect -6 -87394 1146 -87218
rect 2 -88934 1440 -88536
rect -4 -89468 1434 -89070
rect 18 -89960 1478 -89572
rect -6 -90512 1476 -90132
<< via3 >>
rect 26685 8732 26909 8736
rect 26685 8276 26689 8732
rect 26689 8276 26905 8732
rect 26905 8276 26909 8732
rect 26685 8272 26909 8276
rect 20125 4214 20189 4278
rect 20205 4214 20269 4278
rect -391 6 -387 70
rect -387 6 -327 70
rect -311 6 -247 70
rect -231 6 -167 70
rect -151 6 -87 70
rect -71 6 -7 70
rect 9 6 69 70
rect 69 6 73 70
rect 23448 -180 23512 -116
rect 23528 -180 23592 -116
rect 23608 -180 23672 -116
rect 23688 -180 23752 -116
rect 32850 -182 32914 -118
rect 32930 -182 32994 -118
rect 33010 -182 33074 -118
rect 33090 -182 33154 -118
rect 33384 -349 33448 -285
rect 33464 -349 33528 -285
rect 33544 -349 33608 -285
rect 33624 -349 33688 -285
rect 33704 -349 33768 -285
rect 33784 -349 33848 -285
rect 20123 -625 20267 -481
rect 34037 -768 34421 -464
rect 1059 -1262 1363 -958
rect 31466 -1270 31610 -966
rect 34635 -1277 35019 -973
rect -367 -7504 97 -7500
rect -367 -7640 -363 -7504
rect -363 -7640 93 -7504
rect 93 -7640 97 -7504
rect -367 -7644 97 -7640
rect 32854 -7636 33158 -7252
rect -356 -7838 188 -7834
rect -356 -7974 -352 -7838
rect -352 -7974 184 -7838
rect 184 -7974 188 -7838
rect -356 -7978 188 -7974
rect 33423 -7834 33807 -7830
rect 33423 -8130 33427 -7834
rect 33427 -8130 33803 -7834
rect 33803 -8130 33807 -7834
rect 33423 -8134 33807 -8130
rect 32433 -10343 32577 -10243
rect 32433 -10467 32437 -10343
rect 32437 -10467 32573 -10343
rect 32573 -10467 32577 -10343
rect -356 -14369 -52 -14225
rect 32238 -14331 32302 -14267
rect 32318 -14331 32382 -14267
rect 32398 -14331 32462 -14267
rect 32478 -14331 32542 -14267
rect 32558 -14331 32622 -14267
rect 32849 -15760 33153 -15296
rect 33412 -16543 33796 -16079
rect 34059 -17365 34443 -16901
rect 34634 -18168 35018 -17704
<< metal4 >>
rect 26684 8736 26910 8770
rect 26684 8272 26685 8736
rect 26909 8272 26910 8736
rect 26684 8238 26910 8272
rect 20094 4278 20302 4318
rect 20094 4214 20125 4278
rect 20189 4214 20205 4278
rect 20269 4214 20302 4278
rect 20094 4166 20302 4214
rect -422 70 112 122
rect -422 6 -391 70
rect -327 6 -311 70
rect -247 6 -231 70
rect -167 6 -151 70
rect -87 6 -71 70
rect -7 6 9 70
rect 73 6 112 70
rect -422 -40 112 6
rect -418 -6709 -218 -40
rect 20094 -481 20300 4166
rect 23440 -116 23760 7980
rect 23440 -180 23448 -116
rect 23512 -180 23528 -116
rect 23592 -180 23608 -116
rect 23672 -180 23688 -116
rect 23752 -180 23760 -116
rect 23440 -194 23760 -180
rect 32806 -118 33202 -104
rect 32806 -182 32850 -118
rect 32914 -182 32930 -118
rect 32994 -182 33010 -118
rect 33074 -182 33090 -118
rect 33154 -182 33202 -118
rect 20094 -625 20123 -481
rect 20267 -625 20300 -481
rect 992 -958 1416 -918
rect 992 -1262 1059 -958
rect 1363 -1262 1416 -958
rect 992 -1613 1416 -1262
rect 992 -1886 1418 -1613
rect 998 -2243 1418 -1886
rect 20094 -2815 20300 -625
rect 31417 -966 31651 -919
rect 31417 -1270 31466 -966
rect 31610 -1270 31651 -966
rect 31417 -2835 31651 -1270
rect -434 -7135 -218 -6709
rect -418 -7469 -218 -7135
rect 32806 -7180 33202 -182
rect 33378 -285 33856 -95
rect 33378 -349 33384 -285
rect 33448 -349 33464 -285
rect 33528 -349 33544 -285
rect 33608 -349 33624 -285
rect 33688 -349 33704 -285
rect 33768 -349 33784 -285
rect 33848 -349 33856 -285
rect 32806 -7252 33218 -7180
rect -420 -7500 164 -7469
rect -420 -7644 -367 -7500
rect 97 -7644 164 -7500
rect -420 -7667 164 -7644
rect 32806 -7636 32854 -7252
rect 33158 -7636 33218 -7252
rect -418 -7669 162 -7667
rect -418 -7671 -218 -7669
rect 32806 -7712 33218 -7636
rect -406 -7814 -198 -7808
rect -406 -7834 240 -7814
rect -406 -7978 -356 -7834
rect 188 -7978 240 -7834
rect -406 -7998 240 -7978
rect -406 -14192 -198 -7998
rect 32420 -10243 32600 -10212
rect 32420 -10467 32433 -10243
rect 32577 -10467 32600 -10243
rect 32420 -10510 32600 -10467
rect -408 -14225 6 -14192
rect 32420 -14196 32598 -10510
rect -408 -14369 -356 -14225
rect -52 -14369 6 -14225
rect -408 -14388 6 -14369
rect 32200 -14267 32630 -14196
rect 32200 -14331 32238 -14267
rect 32302 -14331 32318 -14267
rect 32382 -14331 32398 -14267
rect 32462 -14331 32478 -14267
rect 32542 -14331 32558 -14267
rect 32622 -14331 32630 -14267
rect 32200 -14406 32630 -14331
rect 32806 -15296 33202 -7712
rect 32806 -15760 32849 -15296
rect 33153 -15760 33202 -15296
rect 32806 -15846 33202 -15760
rect 33378 -7778 33856 -349
rect 33994 -464 34472 -103
rect 33994 -768 34037 -464
rect 34421 -768 34472 -464
rect 33378 -7830 33860 -7778
rect 33378 -8134 33423 -7830
rect 33807 -8134 33860 -7830
rect 33378 -8190 33860 -8134
rect 33378 -16079 33856 -8190
rect 33378 -16543 33412 -16079
rect 33796 -16543 33856 -16079
rect 33378 -16617 33856 -16543
rect 33994 -16901 34472 -768
rect 33994 -17365 34059 -16901
rect 34443 -17365 34472 -16901
rect 33994 -17415 34472 -17365
rect 34596 -973 35074 -100
rect 34596 -1277 34635 -973
rect 35019 -1277 35074 -973
rect 34596 -17704 35074 -1277
rect 34596 -18168 34634 -17704
rect 35018 -18168 35074 -17704
rect 34596 -18217 35074 -18168
use EF_AMUX0801WISO  EF_AMUX0801WISO_0
timestamp 1699118715
transform 1 0 306 0 -1 11000
box -306 -2006 33704 11044
use EF_DACSCA1001  EF_DACSCA1001_0
timestamp 1699118715
transform 1 0 946 0 1 -83429
box -946 -8732 66618 68998
use EF_R2RVCE  EF_R2RVCE_0
timestamp 1699118715
transform 1 0 20662 0 1 -12605
box -804 -1465 11921 11144
use sample_and_hold  sample_and_hold_0
timestamp 1699118715
transform 1 0 -36 0 1 -12655
box 0 -114 19469 11183
<< labels >>
flabel metal3 s 33702 6816 34010 6876 0 FreeSans 60 0 0 0 B[0]
port 1 nsew
flabel metal3 s 33700 6678 34008 6738 0 FreeSans 60 0 0 0 B[1]
port 2 nsew
flabel metal3 s 33704 6544 34012 6604 0 FreeSans 60 0 0 0 B[2]
port 3 nsew
flabel metal2 s 26752 12698 26843 12996 0 FreeSans 60 0 0 0 VIN[0]
port 4 nsew
flabel metal2 s 23308 12698 23404 13000 0 FreeSans 60 0 0 0 VIN[1]
port 5 nsew
flabel metal2 s 20004 12702 20100 13004 0 FreeSans 60 0 0 0 VIN[2]
port 6 nsew
flabel metal2 s 16628 12706 16720 13002 0 FreeSans 60 0 0 0 VIN[3]
port 7 nsew
flabel metal2 s 13318 12700 13410 12996 0 FreeSans 60 0 0 0 VIN[4]
port 8 nsew
flabel metal2 s 10014 12702 10106 12998 0 FreeSans 60 0 0 0 VIN[5]
port 9 nsew
flabel metal2 s 6616 12702 6708 12998 0 FreeSans 60 0 0 0 VIN[6]
port 10 nsew
flabel metal2 s 3218 12706 3310 13002 0 FreeSans 60 0 0 0 VIN[7]
port 11 nsew
flabel metal3 s -1208 -3746 -578 -3544 0 FreeSans 3906 0 0 0 HOLD
port 12 nsew
flabel metal1 s -36 -3749 164 -3549 0 FreeSans 60 0 0 0 HOLD
port 12 nsew
flabel metal3 s 33588 -8490 34002 -8292 0 FreeSans 235 0 0 0 CMP
port 13 nsew
flabel metal3 s -6 -26596 1146 -26420 0 FreeSans 4883 0 0 0 DATA[9]
port 14 nsew
flabel metal3 s -2 -33322 1150 -33146 0 FreeSans 4883 0 0 0 DATA[8]
port 15 nsew
flabel metal3 s -10 -40038 1142 -39862 0 FreeSans 4883 0 0 0 DATA[7]
port 16 nsew
flabel metal3 s 2 -46732 1154 -46556 0 FreeSans 4883 0 0 0 DATA[6]
port 17 nsew
flabel metal3 s 6 -53502 1158 -53326 0 FreeSans 4883 0 0 0 DATA[5]
port 18 nsew
flabel metal3 s -6 -60488 1146 -60312 0 FreeSans 4883 0 0 0 DATA[0]
port 19 nsew
flabel metal3 s 2 -67194 1154 -67018 0 FreeSans 4883 0 0 0 DATA[1]
port 20 nsew
flabel metal3 s -2 -73914 1150 -73738 0 FreeSans 4883 0 0 0 DATA[2]
port 21 nsew
flabel metal3 s -10 -80616 1142 -80440 0 FreeSans 4883 0 0 0 DATA[3]
port 22 nsew
flabel metal3 s -6 -87394 1146 -87218 0 FreeSans 4883 0 0 0 DATA[4]
port 23 nsew
flabel metal3 s -6 -54414 1146 -54238 0 FreeSans 4883 0 0 0 VH
port 24 nsew
flabel metal3 s -16 -54880 1136 -54704 0 FreeSans 4883 0 0 0 VL
port 25 nsew
flabel metal3 s -406 -15086 414 -14884 0 FreeSans 4883 0 0 0 RST
port 26 nsew
flabel metal3 s 2 -88934 1440 -88536 0 FreeSans 4883 0 0 0 DVDD
port 27 nsew
flabel metal3 s -4 -89468 1434 -89070 0 FreeSans 4883 0 0 0 DVSS
port 28 nsew
flabel metal3 s -6 -90512 1476 -90132 0 FreeSans 3125 0 0 0 VSS
port 29 nsew
flabel metal3 s 18 -89960 1478 -89572 0 FreeSans 3125 0 0 0 VDD
port 30 nsew
flabel metal3 s -1208 -7992 -650 -7806 0 FreeSans 3125 0 0 0 EN
port 31 nsew
<< end >>
