VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO EF_ADCS1008NC
  CLASS BLOCK ;
  FOREIGN EF_ADCS1008NC ;
  ORIGIN 0.000 0.000 ;
  SIZE 343.870 BY 517.625 ;
  PIN HOLD
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT 5.870 433.850 6.870 434.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 433.865 3.200 434.875 ;
    END
  END HOLD
  PIN VIN[0]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 139.810 516.085 140.250 517.625 ;
    END
  END VIN[0]
  PIN VIN[1]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 122.580 516.095 123.060 517.625 ;
    END
  END VIN[1]
  PIN VIN[2]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 106.070 516.095 106.550 517.625 ;
    END
  END VIN[2]
  PIN VIN[3]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 89.200 516.095 89.680 517.625 ;
    END
  END VIN[3]
  PIN VIN[4]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 72.640 516.085 73.090 517.625 ;
    END
  END VIN[4]
  PIN VIN[5]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 56.150 516.085 56.600 517.625 ;
    END
  END VIN[5]
  PIN VIN[6]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 39.140 516.125 39.590 517.625 ;
    END
  END VIN[6]
  PIN VIN[7]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 22.120 516.135 22.600 517.625 ;
    END
  END VIN[7]
  PIN EN
    ANTENNAGATEAREA 1.752000 ;
    ANTENNADIFFAREA 1.080000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.635 2.800 413.565 ;
    END
  END EN
  PIN RST
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.165 2.500 378.175 ;
    END
  END RST
  PIN DATA[9]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.615 2.770 320.495 ;
    END
  END DATA[9]
  PIN DATA[8]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.985 3.240 286.865 ;
    END
  END DATA[8]
  PIN DATA[7]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.405 3.240 253.285 ;
    END
  END DATA[7]
  PIN DATA[6]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.935 3.240 219.815 ;
    END
  END DATA[6]
  PIN DATA[5]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.085 3.240 185.965 ;
    END
  END DATA[5]
  PIN DATA[0]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.155 3.240 151.035 ;
    END
  END DATA[0]
  PIN DATA[1]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.625 3.240 117.505 ;
    END
  END DATA[1]
  PIN DATA[2]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.025 3.240 83.905 ;
    END
  END DATA[2]
  PIN DATA[3]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.515 3.240 50.395 ;
    END
  END DATA[3]
  PIN DATA[4]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.625 3.240 16.505 ;
    END
  END DATA[4]
  PIN DVSS
    ANTENNAGATEAREA 74.759102 ;
    ANTENNADIFFAREA 1023.766663 ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.255 4.440 7.255 ;
    END
  END DVSS
  PIN DVDD
    ANTENNAGATEAREA 47.261497 ;
    ANTENNADIFFAREA 93.596451 ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.935 4.440 9.935 ;
    END
  END DVDD
  PIN VDD
    ANTENNAGATEAREA 100.000000 ;
    ANTENNADIFFAREA 2509.495605 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.795 4.620 4.755 ;
    END
  END VDD
  PIN VH
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.525 3.290 181.405 ;
    END
  END VH
  PIN VL
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.195 3.290 179.075 ;
    END
  END VL
  PIN B[0]
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 175.980 516.705 176.280 517.625 ;
    END
  END B[0]
  PIN B[1]
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 176.710 516.685 177.010 517.625 ;
    END
  END B[1]
  PIN B[2]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 177.440 516.685 177.740 517.625 ;
    END
  END B[2]
  PIN CMP
    ANTENNADIFFAREA 0.492900 ;
    PORT
      LAYER met2 ;
        RECT 182.020 515.425 182.990 517.625 ;
    END
  END CMP
  PIN VSS
    ANTENNAGATEAREA 130.500000 ;
    ANTENNADIFFAREA 621.362671 ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.000 6.120 1.930 ;
    END
  END VSS
  OBS
      LAYER li1 ;
        RECT 7.235 14.075 247.920 507.390 ;
      LAYER met1 ;
        RECT 0.055 435.130 248.615 507.595 ;
        RECT 0.055 433.570 5.590 435.130 ;
        RECT 7.150 433.570 248.615 435.130 ;
        RECT 0.055 11.760 248.615 433.570 ;
      LAYER met2 ;
        RECT 0.010 515.855 21.840 517.600 ;
        RECT 22.880 515.855 38.860 517.600 ;
        RECT 0.010 515.845 38.860 515.855 ;
        RECT 39.870 515.845 55.870 517.600 ;
        RECT 0.010 515.805 55.870 515.845 ;
        RECT 56.880 515.805 72.360 517.600 ;
        RECT 73.370 515.815 88.920 517.600 ;
        RECT 89.960 515.815 105.790 517.600 ;
        RECT 106.830 515.815 122.300 517.600 ;
        RECT 123.340 515.815 139.530 517.600 ;
        RECT 73.370 515.805 139.530 515.815 ;
        RECT 140.530 516.425 175.700 517.600 ;
        RECT 140.530 516.405 176.430 516.425 ;
        RECT 178.020 516.405 181.740 517.600 ;
        RECT 140.530 515.805 181.740 516.405 ;
        RECT 0.010 515.145 181.740 515.805 ;
        RECT 183.270 515.145 246.300 517.600 ;
        RECT 0.010 11.760 246.300 515.145 ;
      LAYER met3 ;
        RECT 0.000 435.275 343.870 517.475 ;
        RECT 3.600 433.465 343.870 435.275 ;
        RECT 0.000 413.965 343.870 433.465 ;
        RECT 3.200 412.235 343.870 413.965 ;
        RECT 0.000 378.575 343.870 412.235 ;
        RECT 2.900 376.765 343.870 378.575 ;
        RECT 0.000 320.895 343.870 376.765 ;
        RECT 3.170 319.215 343.870 320.895 ;
        RECT 0.000 287.265 343.870 319.215 ;
        RECT 3.640 285.585 343.870 287.265 ;
        RECT 0.000 253.685 343.870 285.585 ;
        RECT 3.640 252.005 343.870 253.685 ;
        RECT 0.000 220.215 343.870 252.005 ;
        RECT 3.640 218.535 343.870 220.215 ;
        RECT 0.000 186.365 343.870 218.535 ;
        RECT 3.640 184.685 343.870 186.365 ;
        RECT 0.000 181.805 343.870 184.685 ;
        RECT 3.690 180.125 343.870 181.805 ;
        RECT 0.000 179.475 343.870 180.125 ;
        RECT 3.690 177.795 343.870 179.475 ;
        RECT 0.000 151.435 343.870 177.795 ;
        RECT 3.640 149.755 343.870 151.435 ;
        RECT 0.000 117.905 343.870 149.755 ;
        RECT 3.640 116.225 343.870 117.905 ;
        RECT 0.000 84.305 343.870 116.225 ;
        RECT 3.640 82.625 343.870 84.305 ;
        RECT 0.000 50.795 343.870 82.625 ;
        RECT 3.640 49.115 343.870 50.795 ;
        RECT 0.000 16.905 343.870 49.115 ;
        RECT 3.640 15.225 343.870 16.905 ;
        RECT 0.000 10.335 343.870 15.225 ;
        RECT 4.840 5.155 343.870 10.335 ;
        RECT 5.020 2.395 343.870 5.155 ;
        RECT 0.000 2.330 343.870 2.395 ;
        RECT 6.520 1.935 343.870 2.330 ;
        RECT 0.000 1.930 343.870 1.935 ;
        RECT 6.520 0.000 343.870 1.930 ;
      LAYER met4 ;
        RECT 3.880 0.000 343.700 515.595 ;
      LAYER met5 ;
        RECT 16.945 384.480 170.975 506.910 ;
  END
END EF_ADCS1008NC
END LIBRARY

