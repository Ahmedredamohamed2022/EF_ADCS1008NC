magic
tech sky130A
magscale 1 2
timestamp 1693827120
<< pwell >>
rect -668 3002 668 3088
rect -668 -3002 -582 3002
rect 582 -3002 668 3002
rect -668 -3088 668 -3002
<< psubdiff >>
rect -642 3028 -527 3062
rect -493 3028 -459 3062
rect -425 3028 -391 3062
rect -357 3028 -323 3062
rect -289 3028 -255 3062
rect -221 3028 -187 3062
rect -153 3028 -119 3062
rect -85 3028 -51 3062
rect -17 3028 17 3062
rect 51 3028 85 3062
rect 119 3028 153 3062
rect 187 3028 221 3062
rect 255 3028 289 3062
rect 323 3028 357 3062
rect 391 3028 425 3062
rect 459 3028 493 3062
rect 527 3028 642 3062
rect -642 2941 -608 3028
rect 608 2941 642 3028
rect -642 2873 -608 2907
rect -642 2805 -608 2839
rect -642 2737 -608 2771
rect -642 2669 -608 2703
rect -642 2601 -608 2635
rect -642 2533 -608 2567
rect -642 2465 -608 2499
rect -642 2397 -608 2431
rect -642 2329 -608 2363
rect -642 2261 -608 2295
rect -642 2193 -608 2227
rect -642 2125 -608 2159
rect -642 2057 -608 2091
rect -642 1989 -608 2023
rect -642 1921 -608 1955
rect -642 1853 -608 1887
rect -642 1785 -608 1819
rect -642 1717 -608 1751
rect -642 1649 -608 1683
rect -642 1581 -608 1615
rect -642 1513 -608 1547
rect -642 1445 -608 1479
rect -642 1377 -608 1411
rect -642 1309 -608 1343
rect -642 1241 -608 1275
rect -642 1173 -608 1207
rect -642 1105 -608 1139
rect -642 1037 -608 1071
rect -642 969 -608 1003
rect -642 901 -608 935
rect -642 833 -608 867
rect -642 765 -608 799
rect -642 697 -608 731
rect -642 629 -608 663
rect -642 561 -608 595
rect -642 493 -608 527
rect -642 425 -608 459
rect -642 357 -608 391
rect -642 289 -608 323
rect -642 221 -608 255
rect -642 153 -608 187
rect -642 85 -608 119
rect -642 17 -608 51
rect -642 -51 -608 -17
rect -642 -119 -608 -85
rect -642 -187 -608 -153
rect -642 -255 -608 -221
rect -642 -323 -608 -289
rect -642 -391 -608 -357
rect -642 -459 -608 -425
rect -642 -527 -608 -493
rect -642 -595 -608 -561
rect -642 -663 -608 -629
rect -642 -731 -608 -697
rect -642 -799 -608 -765
rect -642 -867 -608 -833
rect -642 -935 -608 -901
rect -642 -1003 -608 -969
rect -642 -1071 -608 -1037
rect -642 -1139 -608 -1105
rect -642 -1207 -608 -1173
rect -642 -1275 -608 -1241
rect -642 -1343 -608 -1309
rect -642 -1411 -608 -1377
rect -642 -1479 -608 -1445
rect -642 -1547 -608 -1513
rect -642 -1615 -608 -1581
rect -642 -1683 -608 -1649
rect -642 -1751 -608 -1717
rect -642 -1819 -608 -1785
rect -642 -1887 -608 -1853
rect -642 -1955 -608 -1921
rect -642 -2023 -608 -1989
rect -642 -2091 -608 -2057
rect -642 -2159 -608 -2125
rect -642 -2227 -608 -2193
rect -642 -2295 -608 -2261
rect -642 -2363 -608 -2329
rect -642 -2431 -608 -2397
rect -642 -2499 -608 -2465
rect -642 -2567 -608 -2533
rect -642 -2635 -608 -2601
rect -642 -2703 -608 -2669
rect -642 -2771 -608 -2737
rect -642 -2839 -608 -2805
rect -642 -2907 -608 -2873
rect 608 2873 642 2907
rect 608 2805 642 2839
rect 608 2737 642 2771
rect 608 2669 642 2703
rect 608 2601 642 2635
rect 608 2533 642 2567
rect 608 2465 642 2499
rect 608 2397 642 2431
rect 608 2329 642 2363
rect 608 2261 642 2295
rect 608 2193 642 2227
rect 608 2125 642 2159
rect 608 2057 642 2091
rect 608 1989 642 2023
rect 608 1921 642 1955
rect 608 1853 642 1887
rect 608 1785 642 1819
rect 608 1717 642 1751
rect 608 1649 642 1683
rect 608 1581 642 1615
rect 608 1513 642 1547
rect 608 1445 642 1479
rect 608 1377 642 1411
rect 608 1309 642 1343
rect 608 1241 642 1275
rect 608 1173 642 1207
rect 608 1105 642 1139
rect 608 1037 642 1071
rect 608 969 642 1003
rect 608 901 642 935
rect 608 833 642 867
rect 608 765 642 799
rect 608 697 642 731
rect 608 629 642 663
rect 608 561 642 595
rect 608 493 642 527
rect 608 425 642 459
rect 608 357 642 391
rect 608 289 642 323
rect 608 221 642 255
rect 608 153 642 187
rect 608 85 642 119
rect 608 17 642 51
rect 608 -51 642 -17
rect 608 -119 642 -85
rect 608 -187 642 -153
rect 608 -255 642 -221
rect 608 -323 642 -289
rect 608 -391 642 -357
rect 608 -459 642 -425
rect 608 -527 642 -493
rect 608 -595 642 -561
rect 608 -663 642 -629
rect 608 -731 642 -697
rect 608 -799 642 -765
rect 608 -867 642 -833
rect 608 -935 642 -901
rect 608 -1003 642 -969
rect 608 -1071 642 -1037
rect 608 -1139 642 -1105
rect 608 -1207 642 -1173
rect 608 -1275 642 -1241
rect 608 -1343 642 -1309
rect 608 -1411 642 -1377
rect 608 -1479 642 -1445
rect 608 -1547 642 -1513
rect 608 -1615 642 -1581
rect 608 -1683 642 -1649
rect 608 -1751 642 -1717
rect 608 -1819 642 -1785
rect 608 -1887 642 -1853
rect 608 -1955 642 -1921
rect 608 -2023 642 -1989
rect 608 -2091 642 -2057
rect 608 -2159 642 -2125
rect 608 -2227 642 -2193
rect 608 -2295 642 -2261
rect 608 -2363 642 -2329
rect 608 -2431 642 -2397
rect 608 -2499 642 -2465
rect 608 -2567 642 -2533
rect 608 -2635 642 -2601
rect 608 -2703 642 -2669
rect 608 -2771 642 -2737
rect 608 -2839 642 -2805
rect 608 -2907 642 -2873
rect -642 -3028 -608 -2941
rect 608 -3028 642 -2941
rect -642 -3062 -527 -3028
rect -493 -3062 -459 -3028
rect -425 -3062 -391 -3028
rect -357 -3062 -323 -3028
rect -289 -3062 -255 -3028
rect -221 -3062 -187 -3028
rect -153 -3062 -119 -3028
rect -85 -3062 -51 -3028
rect -17 -3062 17 -3028
rect 51 -3062 85 -3028
rect 119 -3062 153 -3028
rect 187 -3062 221 -3028
rect 255 -3062 289 -3028
rect 323 -3062 357 -3028
rect 391 -3062 425 -3028
rect 459 -3062 493 -3028
rect 527 -3062 642 -3028
<< psubdiffcont >>
rect -527 3028 -493 3062
rect -459 3028 -425 3062
rect -391 3028 -357 3062
rect -323 3028 -289 3062
rect -255 3028 -221 3062
rect -187 3028 -153 3062
rect -119 3028 -85 3062
rect -51 3028 -17 3062
rect 17 3028 51 3062
rect 85 3028 119 3062
rect 153 3028 187 3062
rect 221 3028 255 3062
rect 289 3028 323 3062
rect 357 3028 391 3062
rect 425 3028 459 3062
rect 493 3028 527 3062
rect -642 2907 -608 2941
rect -642 2839 -608 2873
rect -642 2771 -608 2805
rect -642 2703 -608 2737
rect -642 2635 -608 2669
rect -642 2567 -608 2601
rect -642 2499 -608 2533
rect -642 2431 -608 2465
rect -642 2363 -608 2397
rect -642 2295 -608 2329
rect -642 2227 -608 2261
rect -642 2159 -608 2193
rect -642 2091 -608 2125
rect -642 2023 -608 2057
rect -642 1955 -608 1989
rect -642 1887 -608 1921
rect -642 1819 -608 1853
rect -642 1751 -608 1785
rect -642 1683 -608 1717
rect -642 1615 -608 1649
rect -642 1547 -608 1581
rect -642 1479 -608 1513
rect -642 1411 -608 1445
rect -642 1343 -608 1377
rect -642 1275 -608 1309
rect -642 1207 -608 1241
rect -642 1139 -608 1173
rect -642 1071 -608 1105
rect -642 1003 -608 1037
rect -642 935 -608 969
rect -642 867 -608 901
rect -642 799 -608 833
rect -642 731 -608 765
rect -642 663 -608 697
rect -642 595 -608 629
rect -642 527 -608 561
rect -642 459 -608 493
rect -642 391 -608 425
rect -642 323 -608 357
rect -642 255 -608 289
rect -642 187 -608 221
rect -642 119 -608 153
rect -642 51 -608 85
rect -642 -17 -608 17
rect -642 -85 -608 -51
rect -642 -153 -608 -119
rect -642 -221 -608 -187
rect -642 -289 -608 -255
rect -642 -357 -608 -323
rect -642 -425 -608 -391
rect -642 -493 -608 -459
rect -642 -561 -608 -527
rect -642 -629 -608 -595
rect -642 -697 -608 -663
rect -642 -765 -608 -731
rect -642 -833 -608 -799
rect -642 -901 -608 -867
rect -642 -969 -608 -935
rect -642 -1037 -608 -1003
rect -642 -1105 -608 -1071
rect -642 -1173 -608 -1139
rect -642 -1241 -608 -1207
rect -642 -1309 -608 -1275
rect -642 -1377 -608 -1343
rect -642 -1445 -608 -1411
rect -642 -1513 -608 -1479
rect -642 -1581 -608 -1547
rect -642 -1649 -608 -1615
rect -642 -1717 -608 -1683
rect -642 -1785 -608 -1751
rect -642 -1853 -608 -1819
rect -642 -1921 -608 -1887
rect -642 -1989 -608 -1955
rect -642 -2057 -608 -2023
rect -642 -2125 -608 -2091
rect -642 -2193 -608 -2159
rect -642 -2261 -608 -2227
rect -642 -2329 -608 -2295
rect -642 -2397 -608 -2363
rect -642 -2465 -608 -2431
rect -642 -2533 -608 -2499
rect -642 -2601 -608 -2567
rect -642 -2669 -608 -2635
rect -642 -2737 -608 -2703
rect -642 -2805 -608 -2771
rect -642 -2873 -608 -2839
rect -642 -2941 -608 -2907
rect 608 2907 642 2941
rect 608 2839 642 2873
rect 608 2771 642 2805
rect 608 2703 642 2737
rect 608 2635 642 2669
rect 608 2567 642 2601
rect 608 2499 642 2533
rect 608 2431 642 2465
rect 608 2363 642 2397
rect 608 2295 642 2329
rect 608 2227 642 2261
rect 608 2159 642 2193
rect 608 2091 642 2125
rect 608 2023 642 2057
rect 608 1955 642 1989
rect 608 1887 642 1921
rect 608 1819 642 1853
rect 608 1751 642 1785
rect 608 1683 642 1717
rect 608 1615 642 1649
rect 608 1547 642 1581
rect 608 1479 642 1513
rect 608 1411 642 1445
rect 608 1343 642 1377
rect 608 1275 642 1309
rect 608 1207 642 1241
rect 608 1139 642 1173
rect 608 1071 642 1105
rect 608 1003 642 1037
rect 608 935 642 969
rect 608 867 642 901
rect 608 799 642 833
rect 608 731 642 765
rect 608 663 642 697
rect 608 595 642 629
rect 608 527 642 561
rect 608 459 642 493
rect 608 391 642 425
rect 608 323 642 357
rect 608 255 642 289
rect 608 187 642 221
rect 608 119 642 153
rect 608 51 642 85
rect 608 -17 642 17
rect 608 -85 642 -51
rect 608 -153 642 -119
rect 608 -221 642 -187
rect 608 -289 642 -255
rect 608 -357 642 -323
rect 608 -425 642 -391
rect 608 -493 642 -459
rect 608 -561 642 -527
rect 608 -629 642 -595
rect 608 -697 642 -663
rect 608 -765 642 -731
rect 608 -833 642 -799
rect 608 -901 642 -867
rect 608 -969 642 -935
rect 608 -1037 642 -1003
rect 608 -1105 642 -1071
rect 608 -1173 642 -1139
rect 608 -1241 642 -1207
rect 608 -1309 642 -1275
rect 608 -1377 642 -1343
rect 608 -1445 642 -1411
rect 608 -1513 642 -1479
rect 608 -1581 642 -1547
rect 608 -1649 642 -1615
rect 608 -1717 642 -1683
rect 608 -1785 642 -1751
rect 608 -1853 642 -1819
rect 608 -1921 642 -1887
rect 608 -1989 642 -1955
rect 608 -2057 642 -2023
rect 608 -2125 642 -2091
rect 608 -2193 642 -2159
rect 608 -2261 642 -2227
rect 608 -2329 642 -2295
rect 608 -2397 642 -2363
rect 608 -2465 642 -2431
rect 608 -2533 642 -2499
rect 608 -2601 642 -2567
rect 608 -2669 642 -2635
rect 608 -2737 642 -2703
rect 608 -2805 642 -2771
rect 608 -2873 642 -2839
rect 608 -2941 642 -2907
rect -527 -3062 -493 -3028
rect -459 -3062 -425 -3028
rect -391 -3062 -357 -3028
rect -323 -3062 -289 -3028
rect -255 -3062 -221 -3028
rect -187 -3062 -153 -3028
rect -119 -3062 -85 -3028
rect -51 -3062 -17 -3028
rect 17 -3062 51 -3028
rect 85 -3062 119 -3028
rect 153 -3062 187 -3028
rect 221 -3062 255 -3028
rect 289 -3062 323 -3028
rect 357 -3062 391 -3028
rect 425 -3062 459 -3028
rect 493 -3062 527 -3028
<< xpolycontact >>
rect -512 2500 -442 2932
rect -512 -2932 -442 -2500
rect -194 2500 -124 2932
rect -194 -2932 -124 -2500
rect 124 2500 194 2932
rect 124 -2932 194 -2500
rect 442 2500 512 2932
rect 442 -2932 512 -2500
<< xpolyres >>
rect -512 -2500 -442 2500
rect -194 -2500 -124 2500
rect 124 -2500 194 2500
rect 442 -2500 512 2500
<< locali >>
rect -642 3028 -527 3062
rect -493 3028 -459 3062
rect -425 3028 -391 3062
rect -357 3028 -323 3062
rect -289 3028 -255 3062
rect -221 3028 -187 3062
rect -153 3028 -119 3062
rect -85 3028 -51 3062
rect -17 3028 17 3062
rect 51 3028 85 3062
rect 119 3028 153 3062
rect 187 3028 221 3062
rect 255 3028 289 3062
rect 323 3028 357 3062
rect 391 3028 425 3062
rect 459 3028 493 3062
rect 527 3028 642 3062
rect -642 2941 -608 3028
rect 608 2941 642 3028
rect -642 2873 -608 2907
rect -642 2805 -608 2839
rect -642 2737 -608 2771
rect -642 2669 -608 2703
rect -642 2601 -608 2635
rect -642 2533 -608 2567
rect 608 2873 642 2907
rect 608 2805 642 2839
rect 608 2737 642 2771
rect 608 2669 642 2703
rect 608 2601 642 2635
rect 608 2533 642 2567
rect -642 2465 -608 2499
rect -642 2397 -608 2431
rect -642 2329 -608 2363
rect -642 2261 -608 2295
rect -642 2193 -608 2227
rect -642 2125 -608 2159
rect -642 2057 -608 2091
rect -642 1989 -608 2023
rect -642 1921 -608 1955
rect -642 1853 -608 1887
rect -642 1785 -608 1819
rect -642 1717 -608 1751
rect -642 1649 -608 1683
rect -642 1581 -608 1615
rect -642 1513 -608 1547
rect -642 1445 -608 1479
rect -642 1377 -608 1411
rect -642 1309 -608 1343
rect -642 1241 -608 1275
rect -642 1173 -608 1207
rect -642 1105 -608 1139
rect -642 1037 -608 1071
rect -642 969 -608 1003
rect -642 901 -608 935
rect -642 833 -608 867
rect -642 765 -608 799
rect -642 697 -608 731
rect -642 629 -608 663
rect -642 561 -608 595
rect -642 493 -608 527
rect -642 425 -608 459
rect -642 357 -608 391
rect -642 289 -608 323
rect -642 221 -608 255
rect -642 153 -608 187
rect -642 85 -608 119
rect -642 17 -608 51
rect -642 -51 -608 -17
rect -642 -119 -608 -85
rect -642 -187 -608 -153
rect -642 -255 -608 -221
rect -642 -323 -608 -289
rect -642 -391 -608 -357
rect -642 -459 -608 -425
rect -642 -527 -608 -493
rect -642 -595 -608 -561
rect -642 -663 -608 -629
rect -642 -731 -608 -697
rect -642 -799 -608 -765
rect -642 -867 -608 -833
rect -642 -935 -608 -901
rect -642 -1003 -608 -969
rect -642 -1071 -608 -1037
rect -642 -1139 -608 -1105
rect -642 -1207 -608 -1173
rect -642 -1275 -608 -1241
rect -642 -1343 -608 -1309
rect -642 -1411 -608 -1377
rect -642 -1479 -608 -1445
rect -642 -1547 -608 -1513
rect -642 -1615 -608 -1581
rect -642 -1683 -608 -1649
rect -642 -1751 -608 -1717
rect -642 -1819 -608 -1785
rect -642 -1887 -608 -1853
rect -642 -1955 -608 -1921
rect -642 -2023 -608 -1989
rect -642 -2091 -608 -2057
rect -642 -2159 -608 -2125
rect -642 -2227 -608 -2193
rect -642 -2295 -608 -2261
rect -642 -2363 -608 -2329
rect -642 -2431 -608 -2397
rect -642 -2499 -608 -2465
rect 608 2465 642 2499
rect 608 2397 642 2431
rect 608 2329 642 2363
rect 608 2261 642 2295
rect 608 2193 642 2227
rect 608 2125 642 2159
rect 608 2057 642 2091
rect 608 1989 642 2023
rect 608 1921 642 1955
rect 608 1853 642 1887
rect 608 1785 642 1819
rect 608 1717 642 1751
rect 608 1649 642 1683
rect 608 1581 642 1615
rect 608 1513 642 1547
rect 608 1445 642 1479
rect 608 1377 642 1411
rect 608 1309 642 1343
rect 608 1241 642 1275
rect 608 1173 642 1207
rect 608 1105 642 1139
rect 608 1037 642 1071
rect 608 969 642 1003
rect 608 901 642 935
rect 608 833 642 867
rect 608 765 642 799
rect 608 697 642 731
rect 608 629 642 663
rect 608 561 642 595
rect 608 493 642 527
rect 608 425 642 459
rect 608 357 642 391
rect 608 289 642 323
rect 608 221 642 255
rect 608 153 642 187
rect 608 85 642 119
rect 608 17 642 51
rect 608 -51 642 -17
rect 608 -119 642 -85
rect 608 -187 642 -153
rect 608 -255 642 -221
rect 608 -323 642 -289
rect 608 -391 642 -357
rect 608 -459 642 -425
rect 608 -527 642 -493
rect 608 -595 642 -561
rect 608 -663 642 -629
rect 608 -731 642 -697
rect 608 -799 642 -765
rect 608 -867 642 -833
rect 608 -935 642 -901
rect 608 -1003 642 -969
rect 608 -1071 642 -1037
rect 608 -1139 642 -1105
rect 608 -1207 642 -1173
rect 608 -1275 642 -1241
rect 608 -1343 642 -1309
rect 608 -1411 642 -1377
rect 608 -1479 642 -1445
rect 608 -1547 642 -1513
rect 608 -1615 642 -1581
rect 608 -1683 642 -1649
rect 608 -1751 642 -1717
rect 608 -1819 642 -1785
rect 608 -1887 642 -1853
rect 608 -1955 642 -1921
rect 608 -2023 642 -1989
rect 608 -2091 642 -2057
rect 608 -2159 642 -2125
rect 608 -2227 642 -2193
rect 608 -2295 642 -2261
rect 608 -2363 642 -2329
rect 608 -2431 642 -2397
rect 608 -2499 642 -2465
rect -642 -2567 -608 -2533
rect -642 -2635 -608 -2601
rect -642 -2703 -608 -2669
rect -642 -2771 -608 -2737
rect -642 -2839 -608 -2805
rect -642 -2907 -608 -2873
rect 608 -2567 642 -2533
rect 608 -2635 642 -2601
rect 608 -2703 642 -2669
rect 608 -2771 642 -2737
rect 608 -2839 642 -2805
rect 608 -2907 642 -2873
rect -642 -3028 -608 -2941
rect 608 -3028 642 -2941
rect -642 -3062 -527 -3028
rect -493 -3062 -459 -3028
rect -425 -3062 -391 -3028
rect -357 -3062 -323 -3028
rect -289 -3062 -255 -3028
rect -221 -3062 -187 -3028
rect -153 -3062 -119 -3028
rect -85 -3062 -51 -3028
rect -17 -3062 17 -3028
rect 51 -3062 85 -3028
rect 119 -3062 153 -3028
rect 187 -3062 221 -3028
rect 255 -3062 289 -3028
rect 323 -3062 357 -3028
rect 391 -3062 425 -3028
rect 459 -3062 493 -3028
rect 527 -3062 642 -3028
<< viali >>
rect -494 2878 -460 2912
rect -494 2806 -460 2840
rect -494 2734 -460 2768
rect -494 2662 -460 2696
rect -494 2590 -460 2624
rect -494 2518 -460 2552
rect -176 2878 -142 2912
rect -176 2806 -142 2840
rect -176 2734 -142 2768
rect -176 2662 -142 2696
rect -176 2590 -142 2624
rect -176 2518 -142 2552
rect 142 2878 176 2912
rect 142 2806 176 2840
rect 142 2734 176 2768
rect 142 2662 176 2696
rect 142 2590 176 2624
rect 142 2518 176 2552
rect 460 2878 494 2912
rect 460 2806 494 2840
rect 460 2734 494 2768
rect 460 2662 494 2696
rect 460 2590 494 2624
rect 460 2518 494 2552
rect -494 -2553 -460 -2519
rect -494 -2625 -460 -2591
rect -494 -2697 -460 -2663
rect -494 -2769 -460 -2735
rect -494 -2841 -460 -2807
rect -494 -2913 -460 -2879
rect -176 -2553 -142 -2519
rect -176 -2625 -142 -2591
rect -176 -2697 -142 -2663
rect -176 -2769 -142 -2735
rect -176 -2841 -142 -2807
rect -176 -2913 -142 -2879
rect 142 -2553 176 -2519
rect 142 -2625 176 -2591
rect 142 -2697 176 -2663
rect 142 -2769 176 -2735
rect 142 -2841 176 -2807
rect 142 -2913 176 -2879
rect 460 -2553 494 -2519
rect 460 -2625 494 -2591
rect 460 -2697 494 -2663
rect 460 -2769 494 -2735
rect 460 -2841 494 -2807
rect 460 -2913 494 -2879
<< metal1 >>
rect -502 2912 -452 2926
rect -502 2878 -494 2912
rect -460 2878 -452 2912
rect -502 2840 -452 2878
rect -502 2806 -494 2840
rect -460 2806 -452 2840
rect -502 2768 -452 2806
rect -502 2734 -494 2768
rect -460 2734 -452 2768
rect -502 2696 -452 2734
rect -502 2662 -494 2696
rect -460 2662 -452 2696
rect -502 2624 -452 2662
rect -502 2590 -494 2624
rect -460 2590 -452 2624
rect -502 2552 -452 2590
rect -502 2518 -494 2552
rect -460 2518 -452 2552
rect -502 2505 -452 2518
rect -184 2912 -134 2926
rect -184 2878 -176 2912
rect -142 2878 -134 2912
rect -184 2840 -134 2878
rect -184 2806 -176 2840
rect -142 2806 -134 2840
rect -184 2768 -134 2806
rect -184 2734 -176 2768
rect -142 2734 -134 2768
rect -184 2696 -134 2734
rect -184 2662 -176 2696
rect -142 2662 -134 2696
rect -184 2624 -134 2662
rect -184 2590 -176 2624
rect -142 2590 -134 2624
rect -184 2552 -134 2590
rect -184 2518 -176 2552
rect -142 2518 -134 2552
rect -184 2505 -134 2518
rect 134 2912 184 2926
rect 134 2878 142 2912
rect 176 2878 184 2912
rect 134 2840 184 2878
rect 134 2806 142 2840
rect 176 2806 184 2840
rect 134 2768 184 2806
rect 134 2734 142 2768
rect 176 2734 184 2768
rect 134 2696 184 2734
rect 134 2662 142 2696
rect 176 2662 184 2696
rect 134 2624 184 2662
rect 134 2590 142 2624
rect 176 2590 184 2624
rect 134 2552 184 2590
rect 134 2518 142 2552
rect 176 2518 184 2552
rect 134 2505 184 2518
rect 452 2912 502 2926
rect 452 2878 460 2912
rect 494 2878 502 2912
rect 452 2840 502 2878
rect 452 2806 460 2840
rect 494 2806 502 2840
rect 452 2768 502 2806
rect 452 2734 460 2768
rect 494 2734 502 2768
rect 452 2696 502 2734
rect 452 2662 460 2696
rect 494 2662 502 2696
rect 452 2624 502 2662
rect 452 2590 460 2624
rect 494 2590 502 2624
rect 452 2552 502 2590
rect 452 2518 460 2552
rect 494 2518 502 2552
rect 452 2505 502 2518
rect -502 -2519 -452 -2505
rect -502 -2553 -494 -2519
rect -460 -2553 -452 -2519
rect -502 -2591 -452 -2553
rect -502 -2625 -494 -2591
rect -460 -2625 -452 -2591
rect -502 -2663 -452 -2625
rect -502 -2697 -494 -2663
rect -460 -2697 -452 -2663
rect -502 -2735 -452 -2697
rect -502 -2769 -494 -2735
rect -460 -2769 -452 -2735
rect -502 -2807 -452 -2769
rect -502 -2841 -494 -2807
rect -460 -2841 -452 -2807
rect -502 -2879 -452 -2841
rect -502 -2913 -494 -2879
rect -460 -2913 -452 -2879
rect -502 -2926 -452 -2913
rect -184 -2519 -134 -2505
rect -184 -2553 -176 -2519
rect -142 -2553 -134 -2519
rect -184 -2591 -134 -2553
rect -184 -2625 -176 -2591
rect -142 -2625 -134 -2591
rect -184 -2663 -134 -2625
rect -184 -2697 -176 -2663
rect -142 -2697 -134 -2663
rect -184 -2735 -134 -2697
rect -184 -2769 -176 -2735
rect -142 -2769 -134 -2735
rect -184 -2807 -134 -2769
rect -184 -2841 -176 -2807
rect -142 -2841 -134 -2807
rect -184 -2879 -134 -2841
rect -184 -2913 -176 -2879
rect -142 -2913 -134 -2879
rect -184 -2926 -134 -2913
rect 134 -2519 184 -2505
rect 134 -2553 142 -2519
rect 176 -2553 184 -2519
rect 134 -2591 184 -2553
rect 134 -2625 142 -2591
rect 176 -2625 184 -2591
rect 134 -2663 184 -2625
rect 134 -2697 142 -2663
rect 176 -2697 184 -2663
rect 134 -2735 184 -2697
rect 134 -2769 142 -2735
rect 176 -2769 184 -2735
rect 134 -2807 184 -2769
rect 134 -2841 142 -2807
rect 176 -2841 184 -2807
rect 134 -2879 184 -2841
rect 134 -2913 142 -2879
rect 176 -2913 184 -2879
rect 134 -2926 184 -2913
rect 452 -2519 502 -2505
rect 452 -2553 460 -2519
rect 494 -2553 502 -2519
rect 452 -2591 502 -2553
rect 452 -2625 460 -2591
rect 494 -2625 502 -2591
rect 452 -2663 502 -2625
rect 452 -2697 460 -2663
rect 494 -2697 502 -2663
rect 452 -2735 502 -2697
rect 452 -2769 460 -2735
rect 494 -2769 502 -2735
rect 452 -2807 502 -2769
rect 452 -2841 460 -2807
rect 494 -2841 502 -2807
rect 452 -2879 502 -2841
rect 452 -2913 460 -2879
rect 494 -2913 502 -2879
rect 452 -2926 502 -2913
<< properties >>
string FIXED_BBOX -625 -3045 625 3045
<< end >>
