magic
tech sky130A
magscale 1 2
timestamp 1699926577
<< metal1 >>
rect 924 91839 1458 91865
rect 924 91807 937 91839
rect 920 91723 937 91807
rect 1437 91807 1458 91839
rect 1437 91723 2426 91807
rect 920 91703 2426 91723
rect 1942 88997 2348 89022
rect 1942 88753 1959 88997
rect 2331 88753 2348 88997
rect 1942 88728 2348 88753
rect 147 88194 1504 88199
rect 147 88172 1510 88194
rect 147 88056 173 88172
rect 737 88056 1510 88172
rect 147 87997 1510 88056
rect 1310 87994 1510 87997
rect 1556 85516 1838 85540
rect 1556 85272 1575 85516
rect 1819 85272 1838 85516
rect 1556 85248 1838 85272
rect 3152 85056 3452 85102
rect 3152 84428 3184 85056
rect 3428 84428 3452 85056
rect 3152 84368 3452 84428
rect 926 84229 1510 84274
rect 926 84113 961 84229
rect 1461 84113 1510 84229
rect 926 84076 1510 84113
rect 948 84074 1510 84076
rect 34716 83953 35206 83961
rect 1304 83929 1510 83938
rect 942 83895 1586 83929
rect 942 83779 980 83895
rect 1544 83779 1586 83895
rect 33440 83915 35206 83953
rect 20782 83861 21130 83866
rect 21204 83861 21398 83865
rect 942 83745 1586 83779
rect 20642 83822 21398 83861
rect 1304 83728 1510 83745
rect 20642 83706 21245 83822
rect 21361 83706 21398 83822
rect 20642 83663 21398 83706
rect 20646 83662 20778 83663
rect 33440 83607 34775 83915
rect 35147 83607 35206 83915
rect 33440 83545 35206 83607
<< via1 >>
rect 937 91723 1437 91839
rect 1959 88753 2331 88997
rect 173 88056 737 88172
rect 1575 85272 1819 85516
rect 3184 84428 3428 85056
rect 961 84113 1461 84229
rect 980 83779 1544 83895
rect 21245 83706 21361 83822
rect 34775 83607 35147 83915
<< metal2 >>
rect 4560 104454 4654 104824
rect 7964 104454 8058 104824
rect 11362 104454 11456 104824
rect 14664 104454 14758 104824
rect 17976 104454 18070 104824
rect 21348 104454 21442 104824
rect 24650 104454 24744 104824
rect 28096 104454 28190 104824
rect 35326 104588 35396 104824
rect 35326 104532 35334 104588
rect 35390 104532 35396 104588
rect 35326 104508 35396 104532
rect 35326 104452 35334 104508
rect 35390 104452 35396 104508
rect 35326 104422 35396 104452
rect 35472 104588 35542 104824
rect 35472 104532 35480 104588
rect 35536 104532 35542 104588
rect 35472 104508 35542 104532
rect 35472 104452 35480 104508
rect 35536 104452 35542 104508
rect 35472 104424 35542 104452
rect 35618 104591 35688 104824
rect 36542 104822 36736 104824
rect 35618 104535 35626 104591
rect 35682 104535 35688 104591
rect 35618 104511 35688 104535
rect 35618 104455 35626 104511
rect 35682 104455 35688 104511
rect 35618 104424 35688 104455
rect 36536 104701 36736 104822
rect 36536 104565 36569 104701
rect 36705 104565 36736 104701
rect 36536 104532 36736 104565
rect 36536 104430 36734 104532
rect 28046 100503 28268 100595
rect 28046 100047 28084 100503
rect 28220 100047 28268 100503
rect 924 91849 1458 91865
rect 924 91839 959 91849
rect 1415 91839 1458 91849
rect 924 91723 937 91839
rect 1437 91723 1458 91839
rect 924 91713 959 91723
rect 1415 91713 1458 91723
rect 924 91703 1458 91713
rect 1922 91629 2258 91639
rect 1922 91573 1941 91629
rect 1997 91573 2021 91629
rect 2077 91573 2101 91629
rect 2157 91573 2181 91629
rect 2237 91573 2258 91629
rect 1546 91450 1856 91470
rect 1546 91394 1591 91450
rect 1647 91394 1671 91450
rect 1727 91394 1751 91450
rect 1807 91394 1856 91450
rect 1546 89042 1856 91394
rect 1544 88712 1856 89042
rect 138 88182 768 88211
rect 138 88172 187 88182
rect 723 88172 768 88182
rect 138 88056 173 88172
rect 737 88056 768 88172
rect 138 88046 187 88056
rect 723 88046 768 88056
rect 138 88009 768 88046
rect 1546 85516 1856 88712
rect 1922 89358 2258 91573
rect 28046 91455 28268 100047
rect 28046 91399 28086 91455
rect 28142 91399 28166 91455
rect 28222 91399 28268 91455
rect 28046 91378 28268 91399
rect 3148 91263 3448 91307
rect 3148 90967 3189 91263
rect 3405 90967 3448 91263
rect 1922 89044 2376 89358
rect 1922 88997 2382 89044
rect 1922 88753 1959 88997
rect 2331 88753 2382 88997
rect 1922 88694 2382 88753
rect 1546 85272 1575 85516
rect 1819 85272 1856 85516
rect 1546 85243 1856 85272
rect 3148 85102 3448 90967
rect 3148 85056 3452 85102
rect 3148 84428 3184 85056
rect 3428 84428 3452 85056
rect 3148 84394 3452 84428
rect 3152 84368 3452 84394
rect 926 84239 1510 84274
rect 926 84229 983 84239
rect 1439 84229 1510 84239
rect 926 84113 961 84229
rect 1461 84113 1510 84229
rect 926 84103 983 84113
rect 1439 84103 1510 84113
rect 926 84076 1510 84103
rect 942 83905 1586 83929
rect 942 83895 994 83905
rect 1530 83895 1586 83905
rect 942 83779 980 83895
rect 1544 83779 1586 83895
rect 34716 83915 35206 83961
rect 34716 83909 34775 83915
rect 35147 83909 35206 83915
rect 942 83769 994 83779
rect 1530 83769 1586 83779
rect 942 83745 1586 83769
rect 21204 83832 21398 83865
rect 21204 83696 21235 83832
rect 21371 83696 21398 83832
rect 21204 83665 21398 83696
rect 34716 83613 34773 83909
rect 35149 83613 35206 83909
rect 34716 83607 34775 83613
rect 35147 83607 35206 83613
rect 34716 83553 35206 83607
rect 33766 81400 33942 81529
rect 33766 81264 33783 81400
rect 33919 81264 33942 81400
rect 33766 81233 33942 81264
rect 19338 78452 19950 78537
rect 19338 77996 19441 78452
rect 19817 77996 19950 78452
rect 19338 77927 19950 77996
rect 19482 77003 19746 77927
rect 23730 77495 24346 77563
rect 23730 77039 23795 77495
rect 24251 77039 24346 77495
rect 32336 77209 32888 77211
rect 19510 76675 19732 77003
rect 23730 76969 24346 77039
rect 32334 77120 32898 77209
rect 23906 76683 24122 76969
rect 32334 76744 32388 77120
rect 32844 76744 32898 77120
rect 32334 76671 32898 76744
rect 32336 76653 32888 76671
rect 32472 76553 32694 76653
<< via2 >>
rect 35334 104532 35390 104588
rect 35334 104452 35390 104508
rect 35480 104532 35536 104588
rect 35480 104452 35536 104508
rect 35626 104535 35682 104591
rect 35626 104455 35682 104511
rect 36569 104565 36705 104701
rect 28084 100047 28220 100503
rect 959 91839 1415 91849
rect 959 91723 1415 91839
rect 959 91713 1415 91723
rect 1941 91573 1997 91629
rect 2021 91573 2077 91629
rect 2101 91573 2157 91629
rect 2181 91573 2237 91629
rect 1591 91394 1647 91450
rect 1671 91394 1727 91450
rect 1751 91394 1807 91450
rect 187 88172 723 88182
rect 187 88056 723 88172
rect 187 88046 723 88056
rect 28086 91399 28142 91455
rect 28166 91399 28222 91455
rect 3189 90967 3405 91263
rect 983 84229 1439 84239
rect 983 84113 1439 84229
rect 983 84103 1439 84113
rect 994 83895 1530 83905
rect 994 83779 1530 83895
rect 994 83769 1530 83779
rect 21235 83822 21371 83832
rect 21235 83706 21245 83822
rect 21245 83706 21361 83822
rect 21361 83706 21371 83822
rect 21235 83696 21371 83706
rect 34773 83613 34775 83909
rect 34775 83613 35147 83909
rect 35147 83613 35149 83909
rect 33783 81264 33919 81400
rect 19441 77996 19817 78452
rect 23795 77039 24251 77495
rect 32388 76744 32844 77120
<< metal3 >>
rect 36542 104701 36734 104794
rect 35326 104588 35396 104624
rect 35326 104532 35334 104588
rect 35390 104532 35396 104588
rect 35326 104508 35396 104532
rect 35326 104452 35334 104508
rect 35390 104452 35396 104508
rect 35326 104422 35396 104452
rect 35472 104588 35542 104626
rect 35472 104532 35480 104588
rect 35536 104532 35542 104588
rect 35472 104508 35542 104532
rect 35472 104452 35480 104508
rect 35536 104452 35542 104508
rect 35472 104424 35542 104452
rect 35618 104591 35688 104626
rect 35618 104535 35626 104591
rect 35682 104535 35688 104591
rect 35618 104511 35688 104535
rect 35618 104455 35626 104511
rect 35682 104455 35688 104511
rect 35618 104424 35688 104455
rect 36542 104565 36569 104701
rect 36705 104565 36734 104701
rect 28068 100507 28244 100562
rect 28068 100503 28120 100507
rect 28184 100503 28244 100507
rect 28068 100047 28084 100503
rect 28220 100047 28244 100503
rect 28068 100043 28120 100047
rect 28184 100043 28244 100047
rect 28068 99984 28244 100043
rect 35332 98619 35392 104422
rect 34938 98559 35392 98619
rect 35477 98481 35538 104424
rect 35046 98421 35538 98481
rect 35243 98420 35538 98421
rect 35243 98419 35499 98420
rect 35624 98347 35684 104424
rect 34948 98287 35684 98347
rect 21440 96021 21648 96061
rect 21440 95957 21471 96021
rect 21535 95957 21551 96021
rect 21615 95957 21648 96021
rect 21440 95909 21648 95957
rect 924 91849 1458 91865
rect 924 91813 959 91849
rect 1415 91813 1458 91849
rect 924 91749 955 91813
rect 1419 91749 1458 91813
rect 924 91713 959 91749
rect 1415 91713 1458 91749
rect 924 91703 1458 91713
rect 1346 91629 36432 91641
rect 1346 91573 1941 91629
rect 1997 91573 2021 91629
rect 2077 91573 2101 91629
rect 2157 91573 2181 91629
rect 2237 91627 36432 91629
rect 2237 91573 24794 91627
rect 1346 91563 24794 91573
rect 24858 91563 24874 91627
rect 24938 91563 24954 91627
rect 25018 91563 25034 91627
rect 25098 91625 36432 91627
rect 25098 91563 34196 91625
rect 1346 91561 34196 91563
rect 34260 91561 34276 91625
rect 34340 91561 34356 91625
rect 34420 91561 34436 91625
rect 34500 91561 36432 91625
rect 1346 91547 36432 91561
rect 1342 91463 36432 91471
rect 1340 91458 36432 91463
rect 1340 91455 34730 91458
rect 1340 91450 28086 91455
rect 1340 91394 1591 91450
rect 1647 91394 1671 91450
rect 1727 91394 1751 91450
rect 1807 91399 28086 91450
rect 28142 91399 28166 91455
rect 28222 91399 34730 91455
rect 1807 91394 34730 91399
rect 34794 91394 34810 91458
rect 34874 91394 34890 91458
rect 34954 91394 34970 91458
rect 35034 91394 35050 91458
rect 35114 91394 35130 91458
rect 35194 91394 36432 91458
rect 1340 91377 36432 91394
rect 1340 91373 1638 91377
rect 1340 91307 2490 91309
rect 1336 91279 36432 91307
rect 1336 91263 35383 91279
rect 1336 90967 3189 91263
rect 3405 91262 35383 91263
rect 3405 91118 21469 91262
rect 21613 91118 35383 91262
rect 3405 90975 35383 91118
rect 35767 90975 36432 91279
rect 3405 90967 36432 90975
rect 1336 90907 36432 90967
rect 1346 90785 36432 90825
rect 1346 90515 2405 90785
rect 1360 90481 2405 90515
rect 2709 90777 36432 90785
rect 2709 90481 32812 90777
rect 1360 90473 32812 90481
rect 32956 90770 36432 90777
rect 32956 90473 35981 90770
rect 1360 90466 35981 90473
rect 36365 90466 36432 90770
rect 1360 90425 36432 90466
rect 136 88182 776 88199
rect 136 88046 187 88182
rect 723 88046 776 88182
rect 136 87997 776 88046
rect 33746 84491 34558 84547
rect 926 84243 1510 84274
rect 926 84099 979 84243
rect 1443 84099 1510 84243
rect 926 84076 1510 84099
rect 33746 84107 34200 84491
rect 34504 84107 34558 84491
rect 33746 84043 34558 84107
rect 136 83931 696 83937
rect 136 83929 1582 83931
rect 136 83909 1586 83929
rect 136 83765 990 83909
rect 1534 83765 1586 83909
rect 34716 83913 35206 83961
rect 136 83751 1586 83765
rect 942 83745 1586 83751
rect 21204 83832 21396 83881
rect 21204 83696 21235 83832
rect 21371 83696 21396 83832
rect 21204 82169 21396 83696
rect 34716 83609 34769 83913
rect 35153 83609 35206 83913
rect 34716 83553 35206 83609
rect 34934 83447 35348 83451
rect 36542 83447 36734 104565
rect 33140 83255 36734 83447
rect 34934 83253 35348 83255
rect 19338 78452 19950 78537
rect 19338 77996 19441 78452
rect 19817 78335 19950 78452
rect 21206 78335 21398 82068
rect 33766 81500 33942 81529
rect 33766 81276 33779 81500
rect 33923 81276 33942 81500
rect 33766 81264 33783 81276
rect 33919 81264 33942 81276
rect 33766 81233 33942 81264
rect 19817 78143 21398 78335
rect 19817 77996 19950 78143
rect 19338 77927 19950 77996
rect 23730 77551 24346 77563
rect 938 77547 33626 77551
rect 938 77518 33976 77547
rect 938 77374 990 77518
rect 1294 77495 33976 77518
rect 1294 77374 23795 77495
rect 938 77355 23795 77374
rect 942 77351 23795 77355
rect 23730 77039 23795 77351
rect 24251 77476 33976 77495
rect 24251 77412 33584 77476
rect 33648 77412 33664 77476
rect 33728 77412 33744 77476
rect 33808 77412 33824 77476
rect 33888 77412 33904 77476
rect 33968 77412 33976 77476
rect 24251 77351 33976 77412
rect 24251 77039 24346 77351
rect 33546 77337 33976 77351
rect 32336 77209 32888 77211
rect 23730 76969 24346 77039
rect 32334 77120 32898 77209
rect 136 76849 1760 76859
rect 32334 76849 32388 77120
rect 136 76744 32388 76849
rect 32844 76744 32898 77120
rect 136 76671 32898 76744
rect 136 76657 32888 76671
rect 32336 76653 32888 76657
rect 34184 76447 34510 76467
rect 34184 75983 34195 76447
rect 34499 75983 34510 76447
rect 34184 75963 34510 75983
rect 34734 75664 35166 75665
rect 34734 75200 34758 75664
rect 35142 75200 35166 75664
rect 34734 75199 35166 75200
rect 35394 74842 35800 74847
rect 35394 74378 35405 74842
rect 35789 74378 35800 74842
rect 35394 74373 35800 74378
rect 35962 74039 36382 74067
rect 35962 73575 35980 74039
rect 36364 73575 36382 74039
rect 35962 73547 36382 73575
rect 136 65147 2492 65323
rect 136 58421 2496 58597
rect 136 51705 2488 51881
rect 136 45011 2500 45187
rect 136 38241 2504 38417
rect 136 37329 2492 37505
rect 136 36863 2482 37039
rect 136 31255 2492 31431
rect 136 24549 2500 24725
rect 136 17829 2496 18005
rect 136 11127 2488 11303
rect 136 4349 2492 4525
rect 136 3206 1024 3211
rect 1348 3206 2786 3207
rect 136 2811 2786 3206
rect 1348 2809 2786 2811
rect 136 2673 1024 2675
rect 136 2275 2780 2673
rect 136 2171 1060 2175
rect 136 1783 2824 2171
rect 136 1600 2822 1611
rect 136 1224 3408 1600
<< via3 >>
rect 28120 100503 28184 100507
rect 28120 100443 28184 100503
rect 28120 100363 28184 100427
rect 28120 100283 28184 100347
rect 28120 100203 28184 100267
rect 28120 100123 28184 100187
rect 28120 100047 28184 100107
rect 28120 100043 28184 100047
rect 21471 95957 21535 96021
rect 21551 95957 21615 96021
rect 955 91749 959 91813
rect 959 91749 1019 91813
rect 1035 91749 1099 91813
rect 1115 91749 1179 91813
rect 1195 91749 1259 91813
rect 1275 91749 1339 91813
rect 1355 91749 1415 91813
rect 1415 91749 1419 91813
rect 24794 91563 24858 91627
rect 24874 91563 24938 91627
rect 24954 91563 25018 91627
rect 25034 91563 25098 91627
rect 34196 91561 34260 91625
rect 34276 91561 34340 91625
rect 34356 91561 34420 91625
rect 34436 91561 34500 91625
rect 34730 91394 34794 91458
rect 34810 91394 34874 91458
rect 34890 91394 34954 91458
rect 34970 91394 35034 91458
rect 35050 91394 35114 91458
rect 35130 91394 35194 91458
rect 21469 91118 21613 91262
rect 35383 90975 35767 91279
rect 2405 90481 2709 90785
rect 32812 90473 32956 90777
rect 35981 90466 36365 90770
rect 979 84239 1443 84243
rect 979 84103 983 84239
rect 983 84103 1439 84239
rect 1439 84103 1443 84239
rect 979 84099 1443 84103
rect 34200 84107 34504 84491
rect 990 83905 1534 83909
rect 990 83769 994 83905
rect 994 83769 1530 83905
rect 1530 83769 1534 83905
rect 990 83765 1534 83769
rect 34769 83909 35153 83913
rect 34769 83613 34773 83909
rect 34773 83613 35149 83909
rect 35149 83613 35153 83909
rect 34769 83609 35153 83613
rect 33779 81400 33923 81500
rect 33779 81276 33783 81400
rect 33783 81276 33919 81400
rect 33919 81276 33923 81400
rect 990 77374 1294 77518
rect 33584 77412 33648 77476
rect 33664 77412 33728 77476
rect 33744 77412 33808 77476
rect 33824 77412 33888 77476
rect 33904 77412 33968 77476
rect 34195 75983 34499 76447
rect 34758 75200 35142 75664
rect 35405 74378 35789 74842
rect 35980 73575 36364 74039
<< metal4 >>
rect 28084 100507 28220 100538
rect 28084 100443 28120 100507
rect 28184 100443 28220 100507
rect 28084 100427 28220 100443
rect 28084 100363 28120 100427
rect 28184 100363 28220 100427
rect 28084 100347 28220 100363
rect 28084 100283 28120 100347
rect 28184 100283 28220 100347
rect 28084 100267 28220 100283
rect 28084 100203 28120 100267
rect 28184 100203 28220 100267
rect 28084 100187 28220 100203
rect 28084 100123 28120 100187
rect 28184 100123 28220 100187
rect 28084 100107 28220 100123
rect 28084 100043 28120 100107
rect 28184 100043 28220 100107
rect 28084 100012 28220 100043
rect 21440 96021 21648 96061
rect 21440 95957 21471 96021
rect 21535 95957 21551 96021
rect 21615 95957 21648 96021
rect 21440 95909 21648 95957
rect 924 91813 1458 91865
rect 924 91749 955 91813
rect 1019 91749 1035 91813
rect 1099 91749 1115 91813
rect 1179 91749 1195 91813
rect 1259 91749 1275 91813
rect 1339 91749 1355 91813
rect 1419 91749 1458 91813
rect 924 91703 1458 91749
rect 928 85034 1128 91703
rect 21440 91262 21646 95909
rect 24786 91627 25106 99688
rect 24786 91563 24794 91627
rect 24858 91563 24874 91627
rect 24938 91563 24954 91627
rect 25018 91563 25034 91627
rect 25098 91563 25106 91627
rect 24786 91549 25106 91563
rect 34152 91625 34548 91639
rect 34152 91561 34196 91625
rect 34260 91561 34276 91625
rect 34340 91561 34356 91625
rect 34420 91561 34436 91625
rect 34500 91561 34548 91625
rect 21440 91118 21469 91262
rect 21613 91118 21646 91262
rect 2338 90785 2762 90825
rect 2338 90481 2405 90785
rect 2709 90481 2762 90785
rect 2338 90130 2762 90481
rect 2338 89857 2764 90130
rect 2344 89500 2764 89857
rect 21440 89948 21646 91118
rect 32763 90777 32997 90824
rect 32763 90473 32812 90777
rect 32956 90473 32997 90777
rect 21440 89032 21768 89948
rect 21440 88928 21646 89032
rect 32763 88908 32997 90473
rect 912 84608 1128 85034
rect 928 84274 1128 84608
rect 34152 84563 34548 91561
rect 34724 91458 35202 91648
rect 34724 91394 34730 91458
rect 34794 91394 34810 91458
rect 34874 91394 34890 91458
rect 34954 91394 34970 91458
rect 35034 91394 35050 91458
rect 35114 91394 35130 91458
rect 35194 91394 35202 91458
rect 34152 84491 34564 84563
rect 926 84243 1510 84274
rect 926 84099 979 84243
rect 1443 84099 1510 84243
rect 926 84076 1510 84099
rect 34152 84107 34200 84491
rect 34504 84107 34564 84491
rect 928 84074 1508 84076
rect 928 84072 1128 84074
rect 34152 84031 34564 84107
rect 940 83929 1148 83935
rect 940 83909 1586 83929
rect 940 83765 990 83909
rect 1534 83765 1586 83909
rect 940 83745 1586 83765
rect 940 77551 1148 83745
rect 33766 81500 33946 81531
rect 33766 81276 33779 81500
rect 33923 81276 33946 81500
rect 33766 81233 33946 81276
rect 938 77518 1352 77551
rect 33766 77547 33944 81233
rect 938 77374 990 77518
rect 1294 77374 1352 77518
rect 938 77355 1352 77374
rect 33546 77476 33976 77547
rect 33546 77412 33584 77476
rect 33648 77412 33664 77476
rect 33728 77412 33744 77476
rect 33808 77412 33824 77476
rect 33888 77412 33904 77476
rect 33968 77412 33976 77476
rect 33546 77337 33976 77412
rect 34152 76447 34548 84031
rect 34152 75983 34195 76447
rect 34499 75983 34548 76447
rect 34152 75897 34548 75983
rect 34724 83965 35202 91394
rect 35340 91279 35818 91640
rect 35340 90975 35383 91279
rect 35767 90975 35818 91279
rect 34724 83913 35206 83965
rect 34724 83609 34769 83913
rect 35153 83609 35206 83913
rect 34724 83553 35206 83609
rect 34724 75664 35202 83553
rect 34724 75200 34758 75664
rect 35142 75200 35202 75664
rect 34724 75126 35202 75200
rect 35340 74842 35818 90975
rect 35340 74378 35405 74842
rect 35789 74378 35818 74842
rect 35340 74328 35818 74378
rect 35942 90770 36420 91643
rect 35942 90466 35981 90770
rect 36365 90466 36420 90770
rect 35942 74039 36420 90466
rect 35942 73575 35980 74039
rect 36364 73575 36420 74039
rect 35942 73526 36420 73575
use EF_AMUX0801WISO  EF_AMUX0801WISO_1
timestamp 1699926577
transform 1 0 1652 0 -1 102746
box -306 -2006 33704 11044
use EF_DACSCA1001  EF_DACSCA1001_0
timestamp 1699926577
transform 1 0 2290 0 1 8316
box -946 -8316 66618 68998
use EF_R2RVC  EF_R2RVC_0
timestamp 1699926577
transform 1 0 21953 0 1 79135
box -1774 -1465 11921 11144
use sample_and_hold  sample_and_hold_0
timestamp 1699926577
transform 1 0 1218 0 1 79086
box 0 -114 19469 11183
<< labels >>
flabel metal3 s 136 87997 776 88199 0 FreeSans 899 0 0 0 HOLD
port 1 nsew
flabel metal1 s 1310 87994 1510 88194 0 FreeSans 49 0 0 0 HOLD
port 1 nsew
flabel metal3 s 136 83751 696 83937 0 FreeSans 899 0 0 0 EN
port 2 nsew
flabel metal3 s 136 76657 636 76859 0 FreeSans 899 0 0 0 RST
port 3 nsew
flabel metal3 s 136 65147 690 65323 0 FreeSans 899 0 0 0 DATA[9]
port 4 nsew
flabel metal3 s 136 58421 784 58597 0 FreeSans 899 0 0 0 DATA[8]
port 5 nsew
flabel metal3 s 136 51705 784 51881 0 FreeSans 899 0 0 0 DATA[7]
port 6 nsew
flabel metal3 s 136 45011 784 45187 0 FreeSans 899 0 0 0 DATA[6]
port 7 nsew
flabel metal3 s 136 38241 784 38417 0 FreeSans 899 0 0 0 DATA[5]
port 8 nsew
flabel metal3 s 136 31255 784 31431 0 FreeSans 899 0 0 0 DATA[0]
port 9 nsew
flabel metal3 s 136 24549 784 24725 0 FreeSans 899 0 0 0 DATA[1]
port 10 nsew
flabel metal3 s 136 17829 784 18005 0 FreeSans 899 0 0 0 DATA[2]
port 11 nsew
flabel metal3 s 136 11127 784 11303 0 FreeSans 899 0 0 0 DATA[3]
port 12 nsew
flabel metal3 s 136 4349 784 4525 0 FreeSans 899 0 0 0 DATA[4]
port 13 nsew
flabel metal3 s 136 2275 1024 2675 0 FreeSans 899 0 0 0 DVSS
port 14 nsew
flabel metal3 s 136 2811 1024 3211 0 FreeSans 899 0 0 0 DVDD
port 15 nsew
flabel metal3 s 136 1783 1060 2175 0 FreeSans 899 0 0 0 VDD
port 16 nsew
flabel metal3 s 136 37329 794 37505 0 FreeSans 899 0 0 0 VH
port 17 nsew
flabel metal3 s 136 36863 794 37039 0 FreeSans 899 0 0 0 VL
port 18 nsew
flabel metal3 s 136 1224 1360 1610 0 FreeSans 2291 0 0 0 VSS
port 19 nsew
flabel metal2 s 36536 104430 36734 104822 0 FreeSans 500 0 0 0 CMP
port 20 nsew
flabel metal2 s 4560 104454 4654 104824 0 FreeSans 500 0 0 0 VIN[7]
port 21 nsew
flabel metal2 s 7964 104454 8058 104824 0 FreeSans 500 0 0 0 VIN[6]
port 22 nsew
flabel metal2 s 11362 104454 11456 104824 0 FreeSans 500 0 0 0 VIN[5]
port 23 nsew
flabel metal2 s 14664 104454 14758 104824 0 FreeSans 500 0 0 0 VIN[4]
port 24 nsew
flabel metal2 s 17976 104454 18070 104824 0 FreeSans 500 0 0 0 VIN[3]
port 25 nsew
flabel metal2 s 21348 104454 21442 104824 0 FreeSans 500 0 0 0 VIN[2]
port 26 nsew
flabel metal2 s 24650 104454 24744 104824 0 FreeSans 500 0 0 0 VIN[1]
port 27 nsew
flabel metal2 s 28096 104454 28190 104824 0 FreeSans 500 0 0 0 VIN[0]
port 28 nsew
flabel metal2 s 35326 104424 35396 104824 0 FreeSans 500 0 0 0 B[0]
port 29 nsew
flabel metal2 s 35472 104424 35542 104824 0 FreeSans 500 0 0 0 B[1]
port 30 nsew
flabel metal2 s 35618 104424 35688 104824 0 FreeSans 500 0 0 0 B[2]
port 31 nsew
<< end >>
