magic
tech sky130A
magscale 1 2
timestamp 1699926577
<< metal3 >>
rect -2486 992 2486 1040
rect -2486 928 2402 992
rect 2466 928 2486 992
rect -2486 912 2486 928
rect -2486 848 2402 912
rect 2466 848 2486 912
rect -2486 832 2486 848
rect -2486 768 2402 832
rect 2466 768 2486 832
rect -2486 752 2486 768
rect -2486 688 2402 752
rect 2466 688 2486 752
rect -2486 672 2486 688
rect -2486 608 2402 672
rect 2466 608 2486 672
rect -2486 592 2486 608
rect -2486 528 2402 592
rect 2466 528 2486 592
rect -2486 512 2486 528
rect -2486 448 2402 512
rect 2466 448 2486 512
rect -2486 432 2486 448
rect -2486 368 2402 432
rect 2466 368 2486 432
rect -2486 352 2486 368
rect -2486 288 2402 352
rect 2466 288 2486 352
rect -2486 272 2486 288
rect -2486 208 2402 272
rect 2466 208 2486 272
rect -2486 192 2486 208
rect -2486 128 2402 192
rect 2466 128 2486 192
rect -2486 112 2486 128
rect -2486 48 2402 112
rect 2466 48 2486 112
rect -2486 32 2486 48
rect -2486 -32 2402 32
rect 2466 -32 2486 32
rect -2486 -48 2486 -32
rect -2486 -112 2402 -48
rect 2466 -112 2486 -48
rect -2486 -128 2486 -112
rect -2486 -192 2402 -128
rect 2466 -192 2486 -128
rect -2486 -208 2486 -192
rect -2486 -272 2402 -208
rect 2466 -272 2486 -208
rect -2486 -288 2486 -272
rect -2486 -352 2402 -288
rect 2466 -352 2486 -288
rect -2486 -368 2486 -352
rect -2486 -432 2402 -368
rect 2466 -432 2486 -368
rect -2486 -448 2486 -432
rect -2486 -512 2402 -448
rect 2466 -512 2486 -448
rect -2486 -528 2486 -512
rect -2486 -592 2402 -528
rect 2466 -592 2486 -528
rect -2486 -608 2486 -592
rect -2486 -672 2402 -608
rect 2466 -672 2486 -608
rect -2486 -688 2486 -672
rect -2486 -752 2402 -688
rect 2466 -752 2486 -688
rect -2486 -768 2486 -752
rect -2486 -832 2402 -768
rect 2466 -832 2486 -768
rect -2486 -848 2486 -832
rect -2486 -912 2402 -848
rect 2466 -912 2486 -848
rect -2486 -928 2486 -912
rect -2486 -992 2402 -928
rect 2466 -992 2486 -928
rect -2486 -1040 2486 -992
<< via3 >>
rect 2402 928 2466 992
rect 2402 848 2466 912
rect 2402 768 2466 832
rect 2402 688 2466 752
rect 2402 608 2466 672
rect 2402 528 2466 592
rect 2402 448 2466 512
rect 2402 368 2466 432
rect 2402 288 2466 352
rect 2402 208 2466 272
rect 2402 128 2466 192
rect 2402 48 2466 112
rect 2402 -32 2466 32
rect 2402 -112 2466 -48
rect 2402 -192 2466 -128
rect 2402 -272 2466 -208
rect 2402 -352 2466 -288
rect 2402 -432 2466 -368
rect 2402 -512 2466 -448
rect 2402 -592 2466 -528
rect 2402 -672 2466 -608
rect 2402 -752 2466 -688
rect 2402 -832 2466 -768
rect 2402 -912 2466 -848
rect 2402 -992 2466 -928
<< mimcap >>
rect -2446 952 2154 1000
rect -2446 -952 -2378 952
rect 2086 -952 2154 952
rect -2446 -1000 2154 -952
<< mimcapcontact >>
rect -2378 -952 2086 952
<< metal4 >>
rect 2386 992 2482 1028
rect -2407 952 2115 961
rect -2407 -952 -2378 952
rect 2086 -952 2115 952
rect -2407 -961 2115 -952
rect 2386 928 2402 992
rect 2466 928 2482 992
rect 2386 912 2482 928
rect 2386 848 2402 912
rect 2466 848 2482 912
rect 2386 832 2482 848
rect 2386 768 2402 832
rect 2466 768 2482 832
rect 2386 752 2482 768
rect 2386 688 2402 752
rect 2466 688 2482 752
rect 2386 672 2482 688
rect 2386 608 2402 672
rect 2466 608 2482 672
rect 2386 592 2482 608
rect 2386 528 2402 592
rect 2466 528 2482 592
rect 2386 512 2482 528
rect 2386 448 2402 512
rect 2466 448 2482 512
rect 2386 432 2482 448
rect 2386 368 2402 432
rect 2466 368 2482 432
rect 2386 352 2482 368
rect 2386 288 2402 352
rect 2466 288 2482 352
rect 2386 272 2482 288
rect 2386 208 2402 272
rect 2466 208 2482 272
rect 2386 192 2482 208
rect 2386 128 2402 192
rect 2466 128 2482 192
rect 2386 112 2482 128
rect 2386 48 2402 112
rect 2466 48 2482 112
rect 2386 32 2482 48
rect 2386 -32 2402 32
rect 2466 -32 2482 32
rect 2386 -48 2482 -32
rect 2386 -112 2402 -48
rect 2466 -112 2482 -48
rect 2386 -128 2482 -112
rect 2386 -192 2402 -128
rect 2466 -192 2482 -128
rect 2386 -208 2482 -192
rect 2386 -272 2402 -208
rect 2466 -272 2482 -208
rect 2386 -288 2482 -272
rect 2386 -352 2402 -288
rect 2466 -352 2482 -288
rect 2386 -368 2482 -352
rect 2386 -432 2402 -368
rect 2466 -432 2482 -368
rect 2386 -448 2482 -432
rect 2386 -512 2402 -448
rect 2466 -512 2482 -448
rect 2386 -528 2482 -512
rect 2386 -592 2402 -528
rect 2466 -592 2482 -528
rect 2386 -608 2482 -592
rect 2386 -672 2402 -608
rect 2466 -672 2482 -608
rect 2386 -688 2482 -672
rect 2386 -752 2402 -688
rect 2466 -752 2482 -688
rect 2386 -768 2482 -752
rect 2386 -832 2402 -768
rect 2466 -832 2482 -768
rect 2386 -848 2482 -832
rect 2386 -912 2402 -848
rect 2466 -912 2482 -848
rect 2386 -928 2482 -912
rect 2386 -992 2402 -928
rect 2466 -992 2482 -928
rect 2386 -1028 2482 -992
<< properties >>
string FIXED_BBOX -2486 -1040 2194 1040
<< end >>
