magic
tech sky130A
magscale 1 2
timestamp 1693827120
<< nwell >>
rect -308 -362 308 362
<< mvpmos >>
rect -50 -64 50 136
<< mvpdiff >>
rect -108 121 -50 136
rect -108 87 -96 121
rect -62 87 -50 121
rect -108 53 -50 87
rect -108 19 -96 53
rect -62 19 -50 53
rect -108 -15 -50 19
rect -108 -49 -96 -15
rect -62 -49 -50 -15
rect -108 -64 -50 -49
rect 50 121 108 136
rect 50 87 62 121
rect 96 87 108 121
rect 50 53 108 87
rect 50 19 62 53
rect 96 19 108 53
rect 50 -15 108 19
rect 50 -49 62 -15
rect 96 -49 108 -15
rect 50 -64 108 -49
<< mvpdiffc >>
rect -96 87 -62 121
rect -96 19 -62 53
rect -96 -49 -62 -15
rect 62 87 96 121
rect 62 19 96 53
rect 62 -49 96 -15
<< mvnsubdiff >>
rect -242 284 242 296
rect -242 250 -119 284
rect -85 250 -51 284
rect -17 250 17 284
rect 51 250 85 284
rect 119 250 242 284
rect -242 238 242 250
rect -242 187 -184 238
rect -242 153 -230 187
rect -196 153 -184 187
rect 184 187 242 238
rect -242 119 -184 153
rect 184 153 196 187
rect 230 153 242 187
rect -242 85 -230 119
rect -196 85 -184 119
rect -242 51 -184 85
rect -242 17 -230 51
rect -196 17 -184 51
rect -242 -17 -184 17
rect -242 -51 -230 -17
rect -196 -51 -184 -17
rect -242 -85 -184 -51
rect 184 119 242 153
rect 184 85 196 119
rect 230 85 242 119
rect 184 51 242 85
rect 184 17 196 51
rect 230 17 242 51
rect 184 -17 242 17
rect 184 -51 196 -17
rect 230 -51 242 -17
rect -242 -119 -230 -85
rect -196 -119 -184 -85
rect -242 -153 -184 -119
rect -242 -187 -230 -153
rect -196 -187 -184 -153
rect 184 -85 242 -51
rect 184 -119 196 -85
rect 230 -119 242 -85
rect 184 -153 242 -119
rect -242 -238 -184 -187
rect 184 -187 196 -153
rect 230 -187 242 -153
rect 184 -238 242 -187
rect -242 -250 242 -238
rect -242 -284 -119 -250
rect -85 -284 -51 -250
rect -17 -284 17 -250
rect 51 -284 85 -250
rect 119 -284 242 -250
rect -242 -296 242 -284
<< mvnsubdiffcont >>
rect -119 250 -85 284
rect -51 250 -17 284
rect 17 250 51 284
rect 85 250 119 284
rect -230 153 -196 187
rect 196 153 230 187
rect -230 85 -196 119
rect -230 17 -196 51
rect -230 -51 -196 -17
rect 196 85 230 119
rect 196 17 230 51
rect 196 -51 230 -17
rect -230 -119 -196 -85
rect -230 -187 -196 -153
rect 196 -119 230 -85
rect 196 -187 230 -153
rect -119 -284 -85 -250
rect -51 -284 -17 -250
rect 17 -284 51 -250
rect 85 -284 119 -250
<< poly >>
rect -50 136 50 162
rect -50 -111 50 -64
rect -50 -145 -17 -111
rect 17 -145 50 -111
rect -50 -161 50 -145
<< polycont >>
rect -17 -145 17 -111
<< locali >>
rect -230 250 -119 284
rect -85 250 -51 284
rect -17 250 17 284
rect 51 250 85 284
rect 119 250 230 284
rect -230 187 -196 250
rect -230 119 -196 153
rect 196 187 230 250
rect -230 51 -196 85
rect -230 -17 -196 17
rect -230 -85 -196 -51
rect -96 121 -62 140
rect -96 53 -62 55
rect -96 17 -62 19
rect -96 -68 -62 -49
rect 62 121 96 140
rect 62 53 96 55
rect 62 17 96 19
rect 62 -68 96 -49
rect 196 119 230 153
rect 196 51 230 85
rect 196 -17 230 17
rect 196 -85 230 -51
rect -230 -153 -196 -119
rect -50 -145 -17 -111
rect 17 -145 50 -111
rect -230 -250 -196 -187
rect 196 -153 230 -119
rect 196 -250 230 -187
rect -230 -284 -119 -250
rect -85 -284 -51 -250
rect -17 -284 17 -250
rect 51 -284 85 -250
rect 119 -284 230 -250
<< viali >>
rect -96 87 -62 89
rect -96 55 -62 87
rect -96 -15 -62 17
rect -96 -17 -62 -15
rect 62 87 96 89
rect 62 55 96 87
rect 62 -15 96 17
rect 62 -17 96 -15
rect -17 -145 17 -111
<< metal1 >>
rect -102 89 -56 136
rect -102 55 -96 89
rect -62 55 -56 89
rect -102 17 -56 55
rect -102 -17 -96 17
rect -62 -17 -56 17
rect -102 -64 -56 -17
rect 56 89 102 136
rect 56 55 62 89
rect 96 55 102 89
rect 56 17 102 55
rect 56 -17 62 17
rect 96 -17 102 17
rect 56 -64 102 -17
rect -46 -111 46 -105
rect -46 -145 -17 -111
rect 17 -145 46 -111
rect -46 -151 46 -145
<< properties >>
string FIXED_BBOX -213 -267 213 267
<< end >>
