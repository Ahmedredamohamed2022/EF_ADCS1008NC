magic
tech sky130A
magscale 1 2
timestamp 1694031861
<< viali >>
rect 1961 6885 1995 6919
rect 489 6817 523 6851
rect 2237 6817 2271 6851
rect 949 6749 983 6783
rect 2053 6273 2087 6307
rect 2237 6205 2271 6239
rect 1133 5729 1167 5763
rect 2053 5729 2087 5763
rect 2421 5661 2455 5695
rect 1317 5525 1351 5559
rect 581 5321 615 5355
rect 765 5321 799 5355
rect 2053 5185 2087 5219
rect 1777 5117 1811 5151
rect 397 5049 431 5083
rect 613 5049 647 5083
rect 1685 4777 1719 4811
rect 2237 4709 2271 4743
rect 949 4641 983 4675
rect 1501 4641 1535 4675
rect 1685 4641 1719 4675
rect 2513 4641 2547 4675
rect 2789 4641 2823 4675
rect 2421 4573 2455 4607
rect 1317 4029 1351 4063
rect 2881 4029 2915 4063
rect 949 3961 983 3995
rect 3065 3893 3099 3927
rect 2237 3689 2271 3723
rect 489 3553 523 3587
rect 1961 3553 1995 3587
rect 2329 3553 2363 3587
rect 2789 3553 2823 3587
rect 1041 3485 1075 3519
rect 1869 3145 1903 3179
rect 1041 3009 1075 3043
rect 1225 2941 1259 2975
rect 2237 2941 2271 2975
rect 1685 2805 1719 2839
rect 1869 2805 1903 2839
rect 1501 2601 1535 2635
rect 2973 2533 3007 2567
rect 673 2465 707 2499
rect 2421 2465 2455 2499
rect 857 2329 891 2363
rect 1869 2329 1903 2363
rect 1317 2261 1351 2295
rect 1501 2261 1535 2295
rect 1133 1853 1167 1887
rect 1593 1853 1627 1887
rect 1961 1853 1995 1887
rect 2789 1853 2823 1887
rect 1225 1717 1259 1751
rect 2973 1717 3007 1751
rect 949 1513 983 1547
rect 1961 1513 1995 1547
rect 1777 1445 1811 1479
rect 3065 1445 3099 1479
rect 765 1377 799 1411
rect 2513 1377 2547 1411
rect 1409 1241 1443 1275
rect 1777 1173 1811 1207
rect 3065 969 3099 1003
rect 673 901 707 935
rect 489 765 523 799
rect 1593 765 1627 799
rect 2881 765 2915 799
rect 2145 697 2179 731
<< metal1 >>
rect 92 7098 3864 7120
rect 92 7046 1210 7098
rect 1262 7046 1274 7098
rect 1326 7046 1338 7098
rect 1390 7046 1402 7098
rect 1454 7046 1466 7098
rect 1518 7046 2482 7098
rect 2534 7046 2546 7098
rect 2598 7046 2610 7098
rect 2662 7046 2674 7098
rect 2726 7046 2738 7098
rect 2790 7046 3864 7098
rect 92 7024 3864 7046
rect 1946 6916 1952 6928
rect 1907 6888 1952 6916
rect 1946 6876 1952 6888
rect 2004 6876 2010 6928
rect 290 6808 296 6860
rect 348 6848 354 6860
rect 477 6851 535 6857
rect 477 6848 489 6851
rect 348 6820 489 6848
rect 348 6808 354 6820
rect 477 6817 489 6820
rect 523 6817 535 6851
rect 2222 6848 2228 6860
rect 2183 6820 2228 6848
rect 477 6811 535 6817
rect 2222 6808 2228 6820
rect 2280 6808 2286 6860
rect 934 6780 940 6792
rect 895 6752 940 6780
rect 934 6740 940 6752
rect 992 6740 998 6792
rect 92 6554 3864 6576
rect 92 6502 574 6554
rect 626 6502 638 6554
rect 690 6502 702 6554
rect 754 6502 766 6554
rect 818 6502 830 6554
rect 882 6502 1846 6554
rect 1898 6502 1910 6554
rect 1962 6502 1974 6554
rect 2026 6502 2038 6554
rect 2090 6502 2102 6554
rect 2154 6502 3118 6554
rect 3170 6502 3182 6554
rect 3234 6502 3246 6554
rect 3298 6502 3310 6554
rect 3362 6502 3374 6554
rect 3426 6502 3864 6554
rect 92 6480 3864 6502
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6304 2099 6307
rect 3510 6304 3516 6316
rect 2087 6276 3516 6304
rect 2087 6273 2099 6276
rect 2041 6267 2099 6273
rect 3510 6264 3516 6276
rect 3568 6264 3574 6316
rect 2225 6239 2283 6245
rect 2225 6205 2237 6239
rect 2271 6236 2283 6239
rect 2314 6236 2320 6248
rect 2271 6208 2320 6236
rect 2271 6205 2283 6208
rect 2225 6199 2283 6205
rect 2314 6196 2320 6208
rect 2372 6196 2378 6248
rect 92 6010 3864 6032
rect 92 5958 1210 6010
rect 1262 5958 1274 6010
rect 1326 5958 1338 6010
rect 1390 5958 1402 6010
rect 1454 5958 1466 6010
rect 1518 5958 2482 6010
rect 2534 5958 2546 6010
rect 2598 5958 2610 6010
rect 2662 5958 2674 6010
rect 2726 5958 2738 6010
rect 2790 5958 3864 6010
rect 92 5936 3864 5958
rect 1118 5760 1124 5772
rect 1079 5732 1124 5760
rect 1118 5720 1124 5732
rect 1176 5720 1182 5772
rect 2041 5763 2099 5769
rect 2041 5729 2053 5763
rect 2087 5729 2099 5763
rect 2041 5723 2099 5729
rect 934 5652 940 5704
rect 992 5692 998 5704
rect 2056 5692 2084 5723
rect 2406 5692 2412 5704
rect 992 5664 2084 5692
rect 2367 5664 2412 5692
rect 992 5652 998 5664
rect 2406 5652 2412 5664
rect 2464 5652 2470 5704
rect 1305 5559 1363 5565
rect 1305 5525 1317 5559
rect 1351 5556 1363 5559
rect 1578 5556 1584 5568
rect 1351 5528 1584 5556
rect 1351 5525 1363 5528
rect 1305 5519 1363 5525
rect 1578 5516 1584 5528
rect 1636 5516 1642 5568
rect 92 5466 3864 5488
rect 92 5414 574 5466
rect 626 5414 638 5466
rect 690 5414 702 5466
rect 754 5414 766 5466
rect 818 5414 830 5466
rect 882 5414 1846 5466
rect 1898 5414 1910 5466
rect 1962 5414 1974 5466
rect 2026 5414 2038 5466
rect 2090 5414 2102 5466
rect 2154 5414 3118 5466
rect 3170 5414 3182 5466
rect 3234 5414 3246 5466
rect 3298 5414 3310 5466
rect 3362 5414 3374 5466
rect 3426 5414 3864 5466
rect 92 5392 3864 5414
rect 569 5355 627 5361
rect 569 5321 581 5355
rect 615 5321 627 5355
rect 569 5315 627 5321
rect 753 5355 811 5361
rect 753 5321 765 5355
rect 799 5352 811 5355
rect 1118 5352 1124 5364
rect 799 5324 1124 5352
rect 799 5321 811 5324
rect 753 5315 811 5321
rect 584 5284 612 5315
rect 1118 5312 1124 5324
rect 1176 5312 1182 5364
rect 1026 5284 1032 5296
rect 584 5256 1032 5284
rect 1026 5244 1032 5256
rect 1084 5244 1090 5296
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5216 2099 5219
rect 3510 5216 3516 5228
rect 2087 5188 3516 5216
rect 2087 5185 2099 5188
rect 2041 5179 2099 5185
rect 3510 5176 3516 5188
rect 3568 5176 3574 5228
rect 1670 5108 1676 5160
rect 1728 5148 1734 5160
rect 1765 5151 1823 5157
rect 1765 5148 1777 5151
rect 1728 5120 1777 5148
rect 1728 5108 1734 5120
rect 1765 5117 1777 5120
rect 1811 5117 1823 5151
rect 1765 5111 1823 5117
rect 385 5083 443 5089
rect 385 5049 397 5083
rect 431 5049 443 5083
rect 385 5043 443 5049
rect 601 5083 659 5089
rect 601 5049 613 5083
rect 647 5080 659 5083
rect 934 5080 940 5092
rect 647 5052 940 5080
rect 647 5049 659 5052
rect 601 5043 659 5049
rect 400 5012 428 5043
rect 934 5040 940 5052
rect 992 5040 998 5092
rect 1762 5012 1768 5024
rect 400 4984 1768 5012
rect 1762 4972 1768 4984
rect 1820 4972 1826 5024
rect 92 4922 3864 4944
rect 92 4870 1210 4922
rect 1262 4870 1274 4922
rect 1326 4870 1338 4922
rect 1390 4870 1402 4922
rect 1454 4870 1466 4922
rect 1518 4870 2482 4922
rect 2534 4870 2546 4922
rect 2598 4870 2610 4922
rect 2662 4870 2674 4922
rect 2726 4870 2738 4922
rect 2790 4870 3864 4922
rect 92 4848 3864 4870
rect 1670 4808 1676 4820
rect 1631 4780 1676 4808
rect 1670 4768 1676 4780
rect 1728 4768 1734 4820
rect 1762 4768 1768 4820
rect 1820 4808 1826 4820
rect 1820 4780 2636 4808
rect 1820 4768 1826 4780
rect 2222 4740 2228 4752
rect 1044 4712 1808 4740
rect 2183 4712 2228 4740
rect 1044 4684 1072 4712
rect 937 4675 995 4681
rect 937 4641 949 4675
rect 983 4672 995 4675
rect 1026 4672 1032 4684
rect 983 4644 1032 4672
rect 983 4641 995 4644
rect 937 4635 995 4641
rect 1026 4632 1032 4644
rect 1084 4632 1090 4684
rect 1489 4675 1547 4681
rect 1489 4641 1501 4675
rect 1535 4641 1547 4675
rect 1670 4672 1676 4684
rect 1631 4644 1676 4672
rect 1489 4635 1547 4641
rect 1504 4604 1532 4635
rect 1670 4632 1676 4644
rect 1728 4632 1734 4684
rect 1780 4672 1808 4712
rect 2222 4700 2228 4712
rect 2280 4700 2286 4752
rect 2501 4675 2559 4681
rect 2501 4672 2513 4675
rect 1780 4644 2513 4672
rect 2501 4641 2513 4644
rect 2547 4641 2559 4675
rect 2608 4672 2636 4780
rect 2777 4675 2835 4681
rect 2777 4672 2789 4675
rect 2608 4644 2789 4672
rect 2501 4635 2559 4641
rect 2777 4641 2789 4644
rect 2823 4672 2835 4675
rect 2958 4672 2964 4684
rect 2823 4644 2964 4672
rect 2823 4641 2835 4644
rect 2777 4635 2835 4641
rect 2958 4632 2964 4644
rect 3016 4632 3022 4684
rect 2222 4604 2228 4616
rect 1504 4576 2228 4604
rect 2222 4564 2228 4576
rect 2280 4604 2286 4616
rect 2406 4604 2412 4616
rect 2280 4576 2412 4604
rect 2280 4564 2286 4576
rect 2406 4564 2412 4576
rect 2464 4564 2470 4616
rect 92 4378 3864 4400
rect 92 4326 574 4378
rect 626 4326 638 4378
rect 690 4326 702 4378
rect 754 4326 766 4378
rect 818 4326 830 4378
rect 882 4326 1846 4378
rect 1898 4326 1910 4378
rect 1962 4326 1974 4378
rect 2026 4326 2038 4378
rect 2090 4326 2102 4378
rect 2154 4326 3118 4378
rect 3170 4326 3182 4378
rect 3234 4326 3246 4378
rect 3298 4326 3310 4378
rect 3362 4326 3374 4378
rect 3426 4326 3864 4378
rect 92 4304 3864 4326
rect 1305 4063 1363 4069
rect 1305 4029 1317 4063
rect 1351 4060 1363 4063
rect 1762 4060 1768 4072
rect 1351 4032 1768 4060
rect 1351 4029 1363 4032
rect 1305 4023 1363 4029
rect 1762 4020 1768 4032
rect 1820 4020 1826 4072
rect 2866 4060 2872 4072
rect 2827 4032 2872 4060
rect 2866 4020 2872 4032
rect 2924 4020 2930 4072
rect 937 3995 995 4001
rect 937 3961 949 3995
rect 983 3992 995 3995
rect 1026 3992 1032 4004
rect 983 3964 1032 3992
rect 983 3961 995 3964
rect 937 3955 995 3961
rect 1026 3952 1032 3964
rect 1084 3952 1090 4004
rect 3053 3927 3111 3933
rect 3053 3893 3065 3927
rect 3099 3924 3111 3927
rect 3510 3924 3516 3936
rect 3099 3896 3516 3924
rect 3099 3893 3111 3896
rect 3053 3887 3111 3893
rect 3510 3884 3516 3896
rect 3568 3884 3574 3936
rect 92 3834 3864 3856
rect 92 3782 1210 3834
rect 1262 3782 1274 3834
rect 1326 3782 1338 3834
rect 1390 3782 1402 3834
rect 1454 3782 1466 3834
rect 1518 3782 2482 3834
rect 2534 3782 2546 3834
rect 2598 3782 2610 3834
rect 2662 3782 2674 3834
rect 2726 3782 2738 3834
rect 2790 3782 3864 3834
rect 92 3760 3864 3782
rect 2225 3723 2283 3729
rect 2225 3689 2237 3723
rect 2271 3720 2283 3723
rect 2314 3720 2320 3732
rect 2271 3692 2320 3720
rect 2271 3689 2283 3692
rect 2225 3683 2283 3689
rect 2314 3680 2320 3692
rect 2372 3680 2378 3732
rect 1026 3612 1032 3664
rect 1084 3652 1090 3664
rect 1084 3624 2360 3652
rect 1084 3612 1090 3624
rect 474 3584 480 3596
rect 435 3556 480 3584
rect 474 3544 480 3556
rect 532 3544 538 3596
rect 1949 3587 2007 3593
rect 1949 3553 1961 3587
rect 1995 3584 2007 3587
rect 2222 3584 2228 3596
rect 1995 3556 2228 3584
rect 1995 3553 2007 3556
rect 1949 3547 2007 3553
rect 2222 3544 2228 3556
rect 2280 3544 2286 3596
rect 2332 3593 2360 3624
rect 2317 3587 2375 3593
rect 2317 3553 2329 3587
rect 2363 3553 2375 3587
rect 2317 3547 2375 3553
rect 2777 3587 2835 3593
rect 2777 3553 2789 3587
rect 2823 3584 2835 3587
rect 2958 3584 2964 3596
rect 2823 3556 2964 3584
rect 2823 3553 2835 3556
rect 2777 3547 2835 3553
rect 2958 3544 2964 3556
rect 3016 3544 3022 3596
rect 1029 3519 1087 3525
rect 1029 3485 1041 3519
rect 1075 3516 1087 3519
rect 1762 3516 1768 3528
rect 1075 3488 1768 3516
rect 1075 3485 1087 3488
rect 1029 3479 1087 3485
rect 1762 3476 1768 3488
rect 1820 3476 1826 3528
rect 92 3290 3864 3312
rect 92 3238 574 3290
rect 626 3238 638 3290
rect 690 3238 702 3290
rect 754 3238 766 3290
rect 818 3238 830 3290
rect 882 3238 1846 3290
rect 1898 3238 1910 3290
rect 1962 3238 1974 3290
rect 2026 3238 2038 3290
rect 2090 3238 2102 3290
rect 2154 3238 3118 3290
rect 3170 3238 3182 3290
rect 3234 3238 3246 3290
rect 3298 3238 3310 3290
rect 3362 3238 3374 3290
rect 3426 3238 3864 3290
rect 92 3216 3864 3238
rect 1857 3179 1915 3185
rect 1857 3145 1869 3179
rect 1903 3176 1915 3179
rect 2314 3176 2320 3188
rect 1903 3148 2320 3176
rect 1903 3145 1915 3148
rect 1857 3139 1915 3145
rect 2314 3136 2320 3148
rect 2372 3136 2378 3188
rect 1029 3043 1087 3049
rect 1029 3009 1041 3043
rect 1075 3040 1087 3043
rect 1394 3040 1400 3052
rect 1075 3012 1400 3040
rect 1075 3009 1087 3012
rect 1029 3003 1087 3009
rect 1394 3000 1400 3012
rect 1452 3000 1458 3052
rect 1118 2932 1124 2984
rect 1176 2972 1182 2984
rect 1213 2975 1271 2981
rect 1213 2972 1225 2975
rect 1176 2944 1225 2972
rect 1176 2932 1182 2944
rect 1213 2941 1225 2944
rect 1259 2941 1271 2975
rect 1213 2935 1271 2941
rect 1762 2932 1768 2984
rect 1820 2972 1826 2984
rect 2225 2975 2283 2981
rect 2225 2972 2237 2975
rect 1820 2944 2237 2972
rect 1820 2932 1826 2944
rect 2225 2941 2237 2944
rect 2271 2941 2283 2975
rect 2225 2935 2283 2941
rect 1670 2836 1676 2848
rect 1631 2808 1676 2836
rect 1670 2796 1676 2808
rect 1728 2796 1734 2848
rect 1854 2836 1860 2848
rect 1815 2808 1860 2836
rect 1854 2796 1860 2808
rect 1912 2796 1918 2848
rect 92 2746 3864 2768
rect 92 2694 1210 2746
rect 1262 2694 1274 2746
rect 1326 2694 1338 2746
rect 1390 2694 1402 2746
rect 1454 2694 1466 2746
rect 1518 2694 2482 2746
rect 2534 2694 2546 2746
rect 2598 2694 2610 2746
rect 2662 2694 2674 2746
rect 2726 2694 2738 2746
rect 2790 2694 3864 2746
rect 92 2672 3864 2694
rect 934 2592 940 2644
rect 992 2632 998 2644
rect 1489 2635 1547 2641
rect 1489 2632 1501 2635
rect 992 2604 1501 2632
rect 992 2592 998 2604
rect 1489 2601 1501 2604
rect 1535 2632 1547 2635
rect 2406 2632 2412 2644
rect 1535 2604 2412 2632
rect 1535 2601 1547 2604
rect 1489 2595 1547 2601
rect 2406 2592 2412 2604
rect 2464 2592 2470 2644
rect 2958 2564 2964 2576
rect 2919 2536 2964 2564
rect 2958 2524 2964 2536
rect 3016 2524 3022 2576
rect 661 2499 719 2505
rect 661 2465 673 2499
rect 707 2496 719 2499
rect 1670 2496 1676 2508
rect 707 2468 1676 2496
rect 707 2465 719 2468
rect 661 2459 719 2465
rect 1670 2456 1676 2468
rect 1728 2456 1734 2508
rect 2409 2499 2467 2505
rect 2409 2496 2421 2499
rect 2240 2468 2421 2496
rect 2240 2372 2268 2468
rect 2409 2465 2421 2468
rect 2455 2465 2467 2499
rect 2409 2459 2467 2465
rect 845 2363 903 2369
rect 845 2329 857 2363
rect 891 2360 903 2363
rect 1670 2360 1676 2372
rect 891 2332 1676 2360
rect 891 2329 903 2332
rect 845 2323 903 2329
rect 1670 2320 1676 2332
rect 1728 2320 1734 2372
rect 1854 2320 1860 2372
rect 1912 2360 1918 2372
rect 2222 2360 2228 2372
rect 1912 2332 2228 2360
rect 1912 2320 1918 2332
rect 2222 2320 2228 2332
rect 2280 2320 2286 2372
rect 934 2252 940 2304
rect 992 2292 998 2304
rect 1305 2295 1363 2301
rect 1305 2292 1317 2295
rect 992 2264 1317 2292
rect 992 2252 998 2264
rect 1305 2261 1317 2264
rect 1351 2261 1363 2295
rect 1305 2255 1363 2261
rect 1489 2295 1547 2301
rect 1489 2261 1501 2295
rect 1535 2292 1547 2295
rect 1762 2292 1768 2304
rect 1535 2264 1768 2292
rect 1535 2261 1547 2264
rect 1489 2255 1547 2261
rect 1762 2252 1768 2264
rect 1820 2252 1826 2304
rect 92 2202 3864 2224
rect 92 2150 574 2202
rect 626 2150 638 2202
rect 690 2150 702 2202
rect 754 2150 766 2202
rect 818 2150 830 2202
rect 882 2150 1846 2202
rect 1898 2150 1910 2202
rect 1962 2150 1974 2202
rect 2026 2150 2038 2202
rect 2090 2150 2102 2202
rect 2154 2150 3118 2202
rect 3170 2150 3182 2202
rect 3234 2150 3246 2202
rect 3298 2150 3310 2202
rect 3362 2150 3374 2202
rect 3426 2150 3864 2202
rect 92 2128 3864 2150
rect 1854 1980 1860 2032
rect 1912 2020 1918 2032
rect 2866 2020 2872 2032
rect 1912 1992 2872 2020
rect 1912 1980 1918 1992
rect 2866 1980 2872 1992
rect 2924 1980 2930 2032
rect 2314 1952 2320 1964
rect 1596 1924 2320 1952
rect 1026 1844 1032 1896
rect 1084 1884 1090 1896
rect 1596 1893 1624 1924
rect 2314 1912 2320 1924
rect 2372 1912 2378 1964
rect 1121 1887 1179 1893
rect 1121 1884 1133 1887
rect 1084 1856 1133 1884
rect 1084 1844 1090 1856
rect 1121 1853 1133 1856
rect 1167 1853 1179 1887
rect 1121 1847 1179 1853
rect 1581 1887 1639 1893
rect 1581 1853 1593 1887
rect 1627 1853 1639 1887
rect 1581 1847 1639 1853
rect 1949 1887 2007 1893
rect 1949 1853 1961 1887
rect 1995 1853 2007 1887
rect 1949 1847 2007 1853
rect 1964 1816 1992 1847
rect 2038 1844 2044 1896
rect 2096 1884 2102 1896
rect 2777 1887 2835 1893
rect 2777 1884 2789 1887
rect 2096 1856 2789 1884
rect 2096 1844 2102 1856
rect 2777 1853 2789 1856
rect 2823 1853 2835 1887
rect 2777 1847 2835 1853
rect 2958 1844 2964 1896
rect 3016 1844 3022 1896
rect 2976 1816 3004 1844
rect 1964 1788 3004 1816
rect 1118 1708 1124 1760
rect 1176 1748 1182 1760
rect 1213 1751 1271 1757
rect 1213 1748 1225 1751
rect 1176 1720 1225 1748
rect 1176 1708 1182 1720
rect 1213 1717 1225 1720
rect 1259 1717 1271 1751
rect 1213 1711 1271 1717
rect 2866 1708 2872 1760
rect 2924 1748 2930 1760
rect 2961 1751 3019 1757
rect 2961 1748 2973 1751
rect 2924 1720 2973 1748
rect 2924 1708 2930 1720
rect 2961 1717 2973 1720
rect 3007 1717 3019 1751
rect 2961 1711 3019 1717
rect 92 1658 3864 1680
rect 92 1606 1210 1658
rect 1262 1606 1274 1658
rect 1326 1606 1338 1658
rect 1390 1606 1402 1658
rect 1454 1606 1466 1658
rect 1518 1606 2482 1658
rect 2534 1606 2546 1658
rect 2598 1606 2610 1658
rect 2662 1606 2674 1658
rect 2726 1606 2738 1658
rect 2790 1606 3864 1658
rect 92 1584 3864 1606
rect 937 1547 995 1553
rect 937 1513 949 1547
rect 983 1544 995 1547
rect 1854 1544 1860 1556
rect 983 1516 1860 1544
rect 983 1513 995 1516
rect 937 1507 995 1513
rect 1854 1504 1860 1516
rect 1912 1504 1918 1556
rect 1949 1547 2007 1553
rect 1949 1513 1961 1547
rect 1995 1544 2007 1547
rect 2038 1544 2044 1556
rect 1995 1516 2044 1544
rect 1995 1513 2007 1516
rect 1949 1507 2007 1513
rect 2038 1504 2044 1516
rect 2096 1504 2102 1556
rect 1486 1436 1492 1488
rect 1544 1476 1550 1488
rect 1765 1479 1823 1485
rect 1765 1476 1777 1479
rect 1544 1448 1777 1476
rect 1544 1436 1550 1448
rect 1765 1445 1777 1448
rect 1811 1476 1823 1479
rect 2222 1476 2228 1488
rect 1811 1448 2228 1476
rect 1811 1445 1823 1448
rect 1765 1439 1823 1445
rect 2222 1436 2228 1448
rect 2280 1436 2286 1488
rect 3053 1479 3111 1485
rect 3053 1445 3065 1479
rect 3099 1476 3111 1479
rect 3602 1476 3608 1488
rect 3099 1448 3608 1476
rect 3099 1445 3111 1448
rect 3053 1439 3111 1445
rect 3602 1436 3608 1448
rect 3660 1436 3666 1488
rect 753 1411 811 1417
rect 753 1377 765 1411
rect 799 1408 811 1411
rect 934 1408 940 1420
rect 799 1380 940 1408
rect 799 1377 811 1380
rect 753 1371 811 1377
rect 934 1368 940 1380
rect 992 1368 998 1420
rect 1670 1368 1676 1420
rect 1728 1408 1734 1420
rect 2501 1411 2559 1417
rect 2501 1408 2513 1411
rect 1728 1380 2513 1408
rect 1728 1368 1734 1380
rect 2501 1377 2513 1380
rect 2547 1377 2559 1411
rect 2501 1371 2559 1377
rect 1397 1275 1455 1281
rect 1397 1241 1409 1275
rect 1443 1272 1455 1275
rect 2406 1272 2412 1284
rect 1443 1244 2412 1272
rect 1443 1241 1455 1244
rect 1397 1235 1455 1241
rect 2406 1232 2412 1244
rect 2464 1232 2470 1284
rect 1762 1204 1768 1216
rect 1723 1176 1768 1204
rect 1762 1164 1768 1176
rect 1820 1164 1826 1216
rect 92 1114 3864 1136
rect 92 1062 574 1114
rect 626 1062 638 1114
rect 690 1062 702 1114
rect 754 1062 766 1114
rect 818 1062 830 1114
rect 882 1062 1846 1114
rect 1898 1062 1910 1114
rect 1962 1062 1974 1114
rect 2026 1062 2038 1114
rect 2090 1062 2102 1114
rect 2154 1062 3118 1114
rect 3170 1062 3182 1114
rect 3234 1062 3246 1114
rect 3298 1062 3310 1114
rect 3362 1062 3374 1114
rect 3426 1062 3864 1114
rect 92 1040 3864 1062
rect 3053 1003 3111 1009
rect 3053 969 3065 1003
rect 3099 1000 3111 1003
rect 3510 1000 3516 1012
rect 3099 972 3516 1000
rect 3099 969 3111 972
rect 3053 963 3111 969
rect 3510 960 3516 972
rect 3568 960 3574 1012
rect 661 935 719 941
rect 661 901 673 935
rect 707 932 719 935
rect 1486 932 1492 944
rect 707 904 1492 932
rect 707 901 719 904
rect 661 895 719 901
rect 1486 892 1492 904
rect 1544 892 1550 944
rect 474 796 480 808
rect 435 768 480 796
rect 474 756 480 768
rect 532 756 538 808
rect 1578 796 1584 808
rect 1539 768 1584 796
rect 1578 756 1584 768
rect 1636 756 1642 808
rect 2866 796 2872 808
rect 2827 768 2872 796
rect 2866 756 2872 768
rect 2924 756 2930 808
rect 2133 731 2191 737
rect 2133 697 2145 731
rect 2179 728 2191 731
rect 2958 728 2964 740
rect 2179 700 2964 728
rect 2179 697 2191 700
rect 2133 691 2191 697
rect 2958 688 2964 700
rect 3016 688 3022 740
rect 92 570 3864 592
rect 92 518 1210 570
rect 1262 518 1274 570
rect 1326 518 1338 570
rect 1390 518 1402 570
rect 1454 518 1466 570
rect 1518 518 2482 570
rect 2534 518 2546 570
rect 2598 518 2610 570
rect 2662 518 2674 570
rect 2726 518 2738 570
rect 2790 518 3864 570
rect 92 496 3864 518
<< via1 >>
rect 1210 7046 1262 7098
rect 1274 7046 1326 7098
rect 1338 7046 1390 7098
rect 1402 7046 1454 7098
rect 1466 7046 1518 7098
rect 2482 7046 2534 7098
rect 2546 7046 2598 7098
rect 2610 7046 2662 7098
rect 2674 7046 2726 7098
rect 2738 7046 2790 7098
rect 1952 6919 2004 6928
rect 1952 6885 1961 6919
rect 1961 6885 1995 6919
rect 1995 6885 2004 6919
rect 1952 6876 2004 6885
rect 296 6808 348 6860
rect 2228 6851 2280 6860
rect 2228 6817 2237 6851
rect 2237 6817 2271 6851
rect 2271 6817 2280 6851
rect 2228 6808 2280 6817
rect 940 6783 992 6792
rect 940 6749 949 6783
rect 949 6749 983 6783
rect 983 6749 992 6783
rect 940 6740 992 6749
rect 574 6502 626 6554
rect 638 6502 690 6554
rect 702 6502 754 6554
rect 766 6502 818 6554
rect 830 6502 882 6554
rect 1846 6502 1898 6554
rect 1910 6502 1962 6554
rect 1974 6502 2026 6554
rect 2038 6502 2090 6554
rect 2102 6502 2154 6554
rect 3118 6502 3170 6554
rect 3182 6502 3234 6554
rect 3246 6502 3298 6554
rect 3310 6502 3362 6554
rect 3374 6502 3426 6554
rect 3516 6264 3568 6316
rect 2320 6196 2372 6248
rect 1210 5958 1262 6010
rect 1274 5958 1326 6010
rect 1338 5958 1390 6010
rect 1402 5958 1454 6010
rect 1466 5958 1518 6010
rect 2482 5958 2534 6010
rect 2546 5958 2598 6010
rect 2610 5958 2662 6010
rect 2674 5958 2726 6010
rect 2738 5958 2790 6010
rect 1124 5763 1176 5772
rect 1124 5729 1133 5763
rect 1133 5729 1167 5763
rect 1167 5729 1176 5763
rect 1124 5720 1176 5729
rect 940 5652 992 5704
rect 2412 5695 2464 5704
rect 2412 5661 2421 5695
rect 2421 5661 2455 5695
rect 2455 5661 2464 5695
rect 2412 5652 2464 5661
rect 1584 5516 1636 5568
rect 574 5414 626 5466
rect 638 5414 690 5466
rect 702 5414 754 5466
rect 766 5414 818 5466
rect 830 5414 882 5466
rect 1846 5414 1898 5466
rect 1910 5414 1962 5466
rect 1974 5414 2026 5466
rect 2038 5414 2090 5466
rect 2102 5414 2154 5466
rect 3118 5414 3170 5466
rect 3182 5414 3234 5466
rect 3246 5414 3298 5466
rect 3310 5414 3362 5466
rect 3374 5414 3426 5466
rect 1124 5312 1176 5364
rect 1032 5244 1084 5296
rect 3516 5176 3568 5228
rect 1676 5108 1728 5160
rect 940 5040 992 5092
rect 1768 4972 1820 5024
rect 1210 4870 1262 4922
rect 1274 4870 1326 4922
rect 1338 4870 1390 4922
rect 1402 4870 1454 4922
rect 1466 4870 1518 4922
rect 2482 4870 2534 4922
rect 2546 4870 2598 4922
rect 2610 4870 2662 4922
rect 2674 4870 2726 4922
rect 2738 4870 2790 4922
rect 1676 4811 1728 4820
rect 1676 4777 1685 4811
rect 1685 4777 1719 4811
rect 1719 4777 1728 4811
rect 1676 4768 1728 4777
rect 1768 4768 1820 4820
rect 2228 4743 2280 4752
rect 1032 4632 1084 4684
rect 1676 4675 1728 4684
rect 1676 4641 1685 4675
rect 1685 4641 1719 4675
rect 1719 4641 1728 4675
rect 1676 4632 1728 4641
rect 2228 4709 2237 4743
rect 2237 4709 2271 4743
rect 2271 4709 2280 4743
rect 2228 4700 2280 4709
rect 2964 4632 3016 4684
rect 2228 4564 2280 4616
rect 2412 4607 2464 4616
rect 2412 4573 2421 4607
rect 2421 4573 2455 4607
rect 2455 4573 2464 4607
rect 2412 4564 2464 4573
rect 574 4326 626 4378
rect 638 4326 690 4378
rect 702 4326 754 4378
rect 766 4326 818 4378
rect 830 4326 882 4378
rect 1846 4326 1898 4378
rect 1910 4326 1962 4378
rect 1974 4326 2026 4378
rect 2038 4326 2090 4378
rect 2102 4326 2154 4378
rect 3118 4326 3170 4378
rect 3182 4326 3234 4378
rect 3246 4326 3298 4378
rect 3310 4326 3362 4378
rect 3374 4326 3426 4378
rect 1768 4020 1820 4072
rect 2872 4063 2924 4072
rect 2872 4029 2881 4063
rect 2881 4029 2915 4063
rect 2915 4029 2924 4063
rect 2872 4020 2924 4029
rect 1032 3952 1084 4004
rect 3516 3884 3568 3936
rect 1210 3782 1262 3834
rect 1274 3782 1326 3834
rect 1338 3782 1390 3834
rect 1402 3782 1454 3834
rect 1466 3782 1518 3834
rect 2482 3782 2534 3834
rect 2546 3782 2598 3834
rect 2610 3782 2662 3834
rect 2674 3782 2726 3834
rect 2738 3782 2790 3834
rect 2320 3680 2372 3732
rect 1032 3612 1084 3664
rect 480 3587 532 3596
rect 480 3553 489 3587
rect 489 3553 523 3587
rect 523 3553 532 3587
rect 480 3544 532 3553
rect 2228 3544 2280 3596
rect 2964 3544 3016 3596
rect 1768 3476 1820 3528
rect 574 3238 626 3290
rect 638 3238 690 3290
rect 702 3238 754 3290
rect 766 3238 818 3290
rect 830 3238 882 3290
rect 1846 3238 1898 3290
rect 1910 3238 1962 3290
rect 1974 3238 2026 3290
rect 2038 3238 2090 3290
rect 2102 3238 2154 3290
rect 3118 3238 3170 3290
rect 3182 3238 3234 3290
rect 3246 3238 3298 3290
rect 3310 3238 3362 3290
rect 3374 3238 3426 3290
rect 2320 3136 2372 3188
rect 1400 3000 1452 3052
rect 1124 2932 1176 2984
rect 1768 2932 1820 2984
rect 1676 2839 1728 2848
rect 1676 2805 1685 2839
rect 1685 2805 1719 2839
rect 1719 2805 1728 2839
rect 1676 2796 1728 2805
rect 1860 2839 1912 2848
rect 1860 2805 1869 2839
rect 1869 2805 1903 2839
rect 1903 2805 1912 2839
rect 1860 2796 1912 2805
rect 1210 2694 1262 2746
rect 1274 2694 1326 2746
rect 1338 2694 1390 2746
rect 1402 2694 1454 2746
rect 1466 2694 1518 2746
rect 2482 2694 2534 2746
rect 2546 2694 2598 2746
rect 2610 2694 2662 2746
rect 2674 2694 2726 2746
rect 2738 2694 2790 2746
rect 940 2592 992 2644
rect 2412 2592 2464 2644
rect 2964 2567 3016 2576
rect 2964 2533 2973 2567
rect 2973 2533 3007 2567
rect 3007 2533 3016 2567
rect 2964 2524 3016 2533
rect 1676 2456 1728 2508
rect 1676 2320 1728 2372
rect 1860 2363 1912 2372
rect 1860 2329 1869 2363
rect 1869 2329 1903 2363
rect 1903 2329 1912 2363
rect 1860 2320 1912 2329
rect 2228 2320 2280 2372
rect 940 2252 992 2304
rect 1768 2252 1820 2304
rect 574 2150 626 2202
rect 638 2150 690 2202
rect 702 2150 754 2202
rect 766 2150 818 2202
rect 830 2150 882 2202
rect 1846 2150 1898 2202
rect 1910 2150 1962 2202
rect 1974 2150 2026 2202
rect 2038 2150 2090 2202
rect 2102 2150 2154 2202
rect 3118 2150 3170 2202
rect 3182 2150 3234 2202
rect 3246 2150 3298 2202
rect 3310 2150 3362 2202
rect 3374 2150 3426 2202
rect 1860 1980 1912 2032
rect 2872 1980 2924 2032
rect 1032 1844 1084 1896
rect 2320 1912 2372 1964
rect 2044 1844 2096 1896
rect 2964 1844 3016 1896
rect 1124 1708 1176 1760
rect 2872 1708 2924 1760
rect 1210 1606 1262 1658
rect 1274 1606 1326 1658
rect 1338 1606 1390 1658
rect 1402 1606 1454 1658
rect 1466 1606 1518 1658
rect 2482 1606 2534 1658
rect 2546 1606 2598 1658
rect 2610 1606 2662 1658
rect 2674 1606 2726 1658
rect 2738 1606 2790 1658
rect 1860 1504 1912 1556
rect 2044 1504 2096 1556
rect 1492 1436 1544 1488
rect 2228 1436 2280 1488
rect 3608 1436 3660 1488
rect 940 1368 992 1420
rect 1676 1368 1728 1420
rect 2412 1232 2464 1284
rect 1768 1207 1820 1216
rect 1768 1173 1777 1207
rect 1777 1173 1811 1207
rect 1811 1173 1820 1207
rect 1768 1164 1820 1173
rect 574 1062 626 1114
rect 638 1062 690 1114
rect 702 1062 754 1114
rect 766 1062 818 1114
rect 830 1062 882 1114
rect 1846 1062 1898 1114
rect 1910 1062 1962 1114
rect 1974 1062 2026 1114
rect 2038 1062 2090 1114
rect 2102 1062 2154 1114
rect 3118 1062 3170 1114
rect 3182 1062 3234 1114
rect 3246 1062 3298 1114
rect 3310 1062 3362 1114
rect 3374 1062 3426 1114
rect 3516 960 3568 1012
rect 1492 892 1544 944
rect 480 799 532 808
rect 480 765 489 799
rect 489 765 523 799
rect 523 765 532 799
rect 480 756 532 765
rect 1584 799 1636 808
rect 1584 765 1593 799
rect 1593 765 1627 799
rect 1627 765 1636 799
rect 1584 756 1636 765
rect 2872 799 2924 808
rect 2872 765 2881 799
rect 2881 765 2915 799
rect 2915 765 2924 799
rect 2872 756 2924 765
rect 2964 688 3016 740
rect 1210 518 1262 570
rect 1274 518 1326 570
rect 1338 518 1390 570
rect 1402 518 1454 570
rect 1466 518 1518 570
rect 2482 518 2534 570
rect 2546 518 2598 570
rect 2610 518 2662 570
rect 2674 518 2726 570
rect 2738 518 2790 570
<< metal2 >>
rect 1950 7240 2006 7249
rect 1950 7175 2006 7184
rect 1210 7100 1518 7120
rect 1210 7098 1216 7100
rect 1272 7098 1296 7100
rect 1352 7098 1376 7100
rect 1432 7098 1456 7100
rect 1512 7098 1518 7100
rect 1272 7046 1274 7098
rect 1454 7046 1456 7098
rect 1210 7044 1216 7046
rect 1272 7044 1296 7046
rect 1352 7044 1376 7046
rect 1432 7044 1456 7046
rect 1512 7044 1518 7046
rect 1210 7024 1518 7044
rect 1964 6934 1992 7175
rect 2482 7100 2790 7120
rect 2482 7098 2488 7100
rect 2544 7098 2568 7100
rect 2624 7098 2648 7100
rect 2704 7098 2728 7100
rect 2784 7098 2790 7100
rect 2544 7046 2546 7098
rect 2726 7046 2728 7098
rect 2482 7044 2488 7046
rect 2544 7044 2568 7046
rect 2624 7044 2648 7046
rect 2704 7044 2728 7046
rect 2784 7044 2790 7046
rect 2482 7024 2790 7044
rect 1952 6928 2004 6934
rect 1952 6870 2004 6876
rect 296 6860 348 6866
rect 296 6802 348 6808
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 308 6633 336 6802
rect 940 6792 992 6798
rect 940 6734 992 6740
rect 294 6624 350 6633
rect 294 6559 350 6568
rect 574 6556 882 6576
rect 574 6554 580 6556
rect 636 6554 660 6556
rect 716 6554 740 6556
rect 796 6554 820 6556
rect 876 6554 882 6556
rect 636 6502 638 6554
rect 818 6502 820 6554
rect 574 6500 580 6502
rect 636 6500 660 6502
rect 716 6500 740 6502
rect 796 6500 820 6502
rect 876 6500 882 6502
rect 574 6480 882 6500
rect 952 5710 980 6734
rect 1846 6556 2154 6576
rect 1846 6554 1852 6556
rect 1908 6554 1932 6556
rect 1988 6554 2012 6556
rect 2068 6554 2092 6556
rect 2148 6554 2154 6556
rect 1908 6502 1910 6554
rect 2090 6502 2092 6554
rect 1846 6500 1852 6502
rect 1908 6500 1932 6502
rect 1988 6500 2012 6502
rect 2068 6500 2092 6502
rect 2148 6500 2154 6502
rect 1846 6480 2154 6500
rect 1210 6012 1518 6032
rect 1210 6010 1216 6012
rect 1272 6010 1296 6012
rect 1352 6010 1376 6012
rect 1432 6010 1456 6012
rect 1512 6010 1518 6012
rect 1272 5958 1274 6010
rect 1454 5958 1456 6010
rect 1210 5956 1216 5958
rect 1272 5956 1296 5958
rect 1352 5956 1376 5958
rect 1432 5956 1456 5958
rect 1512 5956 1518 5958
rect 1210 5936 1518 5956
rect 1124 5772 1176 5778
rect 1124 5714 1176 5720
rect 940 5704 992 5710
rect 940 5646 992 5652
rect 574 5468 882 5488
rect 574 5466 580 5468
rect 636 5466 660 5468
rect 716 5466 740 5468
rect 796 5466 820 5468
rect 876 5466 882 5468
rect 636 5414 638 5466
rect 818 5414 820 5466
rect 574 5412 580 5414
rect 636 5412 660 5414
rect 716 5412 740 5414
rect 796 5412 820 5414
rect 876 5412 882 5414
rect 574 5392 882 5412
rect 952 5098 980 5646
rect 1136 5370 1164 5714
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 1124 5364 1176 5370
rect 1124 5306 1176 5312
rect 1032 5296 1084 5302
rect 1032 5238 1084 5244
rect 940 5092 992 5098
rect 940 5034 992 5040
rect 574 4380 882 4400
rect 574 4378 580 4380
rect 636 4378 660 4380
rect 716 4378 740 4380
rect 796 4378 820 4380
rect 876 4378 882 4380
rect 636 4326 638 4378
rect 818 4326 820 4378
rect 574 4324 580 4326
rect 636 4324 660 4326
rect 716 4324 740 4326
rect 796 4324 820 4326
rect 876 4324 882 4326
rect 574 4304 882 4324
rect 478 3904 534 3913
rect 478 3839 534 3848
rect 492 3602 520 3839
rect 480 3596 532 3602
rect 480 3538 532 3544
rect 574 3292 882 3312
rect 574 3290 580 3292
rect 636 3290 660 3292
rect 716 3290 740 3292
rect 796 3290 820 3292
rect 876 3290 882 3292
rect 636 3238 638 3290
rect 818 3238 820 3290
rect 574 3236 580 3238
rect 636 3236 660 3238
rect 716 3236 740 3238
rect 796 3236 820 3238
rect 876 3236 882 3238
rect 574 3216 882 3236
rect 952 2650 980 5034
rect 1044 4690 1072 5238
rect 1210 4924 1518 4944
rect 1210 4922 1216 4924
rect 1272 4922 1296 4924
rect 1352 4922 1376 4924
rect 1432 4922 1456 4924
rect 1512 4922 1518 4924
rect 1272 4870 1274 4922
rect 1454 4870 1456 4922
rect 1210 4868 1216 4870
rect 1272 4868 1296 4870
rect 1352 4868 1376 4870
rect 1432 4868 1456 4870
rect 1512 4868 1518 4870
rect 1210 4848 1518 4868
rect 1032 4684 1084 4690
rect 1032 4626 1084 4632
rect 1044 4010 1072 4626
rect 1032 4004 1084 4010
rect 1032 3946 1084 3952
rect 1044 3670 1072 3946
rect 1210 3836 1518 3856
rect 1210 3834 1216 3836
rect 1272 3834 1296 3836
rect 1352 3834 1376 3836
rect 1432 3834 1456 3836
rect 1512 3834 1518 3836
rect 1272 3782 1274 3834
rect 1454 3782 1456 3834
rect 1210 3780 1216 3782
rect 1272 3780 1296 3782
rect 1352 3780 1376 3782
rect 1432 3780 1456 3782
rect 1512 3780 1518 3782
rect 1210 3760 1518 3780
rect 1032 3664 1084 3670
rect 1032 3606 1084 3612
rect 940 2644 992 2650
rect 940 2586 992 2592
rect 940 2304 992 2310
rect 940 2246 992 2252
rect 574 2204 882 2224
rect 574 2202 580 2204
rect 636 2202 660 2204
rect 716 2202 740 2204
rect 796 2202 820 2204
rect 876 2202 882 2204
rect 636 2150 638 2202
rect 818 2150 820 2202
rect 574 2148 580 2150
rect 636 2148 660 2150
rect 716 2148 740 2150
rect 796 2148 820 2150
rect 876 2148 882 2150
rect 574 2128 882 2148
rect 952 1426 980 2246
rect 1044 1902 1072 3606
rect 1398 3496 1454 3505
rect 1398 3431 1454 3440
rect 1412 3058 1440 3431
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1124 2984 1176 2990
rect 1124 2926 1176 2932
rect 1032 1896 1084 1902
rect 1032 1838 1084 1844
rect 1136 1766 1164 2926
rect 1210 2748 1518 2768
rect 1210 2746 1216 2748
rect 1272 2746 1296 2748
rect 1352 2746 1376 2748
rect 1432 2746 1456 2748
rect 1512 2746 1518 2748
rect 1272 2694 1274 2746
rect 1454 2694 1456 2746
rect 1210 2692 1216 2694
rect 1272 2692 1296 2694
rect 1352 2692 1376 2694
rect 1432 2692 1456 2694
rect 1512 2692 1518 2694
rect 1210 2672 1518 2692
rect 1124 1760 1176 1766
rect 1124 1702 1176 1708
rect 1210 1660 1518 1680
rect 1210 1658 1216 1660
rect 1272 1658 1296 1660
rect 1352 1658 1376 1660
rect 1432 1658 1456 1660
rect 1512 1658 1518 1660
rect 1272 1606 1274 1658
rect 1454 1606 1456 1658
rect 1210 1604 1216 1606
rect 1272 1604 1296 1606
rect 1352 1604 1376 1606
rect 1432 1604 1456 1606
rect 1512 1604 1518 1606
rect 1210 1584 1518 1604
rect 1492 1488 1544 1494
rect 1492 1430 1544 1436
rect 940 1420 992 1426
rect 940 1362 992 1368
rect 478 1320 534 1329
rect 478 1255 534 1264
rect 492 814 520 1255
rect 574 1116 882 1136
rect 574 1114 580 1116
rect 636 1114 660 1116
rect 716 1114 740 1116
rect 796 1114 820 1116
rect 876 1114 882 1116
rect 636 1062 638 1114
rect 818 1062 820 1114
rect 574 1060 580 1062
rect 636 1060 660 1062
rect 716 1060 740 1062
rect 796 1060 820 1062
rect 876 1060 882 1062
rect 574 1040 882 1060
rect 1504 950 1532 1430
rect 1492 944 1544 950
rect 1492 886 1544 892
rect 1596 814 1624 5510
rect 1846 5468 2154 5488
rect 1846 5466 1852 5468
rect 1908 5466 1932 5468
rect 1988 5466 2012 5468
rect 2068 5466 2092 5468
rect 2148 5466 2154 5468
rect 1908 5414 1910 5466
rect 2090 5414 2092 5466
rect 1846 5412 1852 5414
rect 1908 5412 1932 5414
rect 1988 5412 2012 5414
rect 2068 5412 2092 5414
rect 2148 5412 2154 5414
rect 1846 5392 2154 5412
rect 1676 5160 1728 5166
rect 1676 5102 1728 5108
rect 1688 4826 1716 5102
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1780 4826 1808 4966
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 1780 4706 1808 4762
rect 2240 4758 2268 6802
rect 3118 6556 3426 6576
rect 3118 6554 3124 6556
rect 3180 6554 3204 6556
rect 3260 6554 3284 6556
rect 3340 6554 3364 6556
rect 3420 6554 3426 6556
rect 3180 6502 3182 6554
rect 3362 6502 3364 6554
rect 3118 6500 3124 6502
rect 3180 6500 3204 6502
rect 3260 6500 3284 6502
rect 3340 6500 3364 6502
rect 3420 6500 3426 6502
rect 3118 6480 3426 6500
rect 3514 6488 3570 6497
rect 3514 6423 3570 6432
rect 3528 6322 3556 6423
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 2320 6248 2372 6254
rect 2320 6190 2372 6196
rect 1688 4690 1808 4706
rect 2228 4752 2280 4758
rect 2228 4694 2280 4700
rect 1676 4684 1808 4690
rect 1728 4678 1808 4684
rect 1676 4626 1728 4632
rect 2228 4616 2280 4622
rect 2228 4558 2280 4564
rect 1846 4380 2154 4400
rect 1846 4378 1852 4380
rect 1908 4378 1932 4380
rect 1988 4378 2012 4380
rect 2068 4378 2092 4380
rect 2148 4378 2154 4380
rect 1908 4326 1910 4378
rect 2090 4326 2092 4378
rect 1846 4324 1852 4326
rect 1908 4324 1932 4326
rect 1988 4324 2012 4326
rect 2068 4324 2092 4326
rect 2148 4324 2154 4326
rect 1846 4304 2154 4324
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1780 3534 1808 4014
rect 2240 3602 2268 4558
rect 2332 3738 2360 6190
rect 2482 6012 2790 6032
rect 2482 6010 2488 6012
rect 2544 6010 2568 6012
rect 2624 6010 2648 6012
rect 2704 6010 2728 6012
rect 2784 6010 2790 6012
rect 2544 5958 2546 6010
rect 2726 5958 2728 6010
rect 2482 5956 2488 5958
rect 2544 5956 2568 5958
rect 2624 5956 2648 5958
rect 2704 5956 2728 5958
rect 2784 5956 2790 5958
rect 2482 5936 2790 5956
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2424 4622 2452 5646
rect 3118 5468 3426 5488
rect 3118 5466 3124 5468
rect 3180 5466 3204 5468
rect 3260 5466 3284 5468
rect 3340 5466 3364 5468
rect 3420 5466 3426 5468
rect 3180 5414 3182 5466
rect 3362 5414 3364 5466
rect 3118 5412 3124 5414
rect 3180 5412 3204 5414
rect 3260 5412 3284 5414
rect 3340 5412 3364 5414
rect 3420 5412 3426 5414
rect 3118 5392 3426 5412
rect 3514 5400 3570 5409
rect 3514 5335 3570 5344
rect 3528 5234 3556 5335
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 2482 4924 2790 4944
rect 2482 4922 2488 4924
rect 2544 4922 2568 4924
rect 2624 4922 2648 4924
rect 2704 4922 2728 4924
rect 2784 4922 2790 4924
rect 2544 4870 2546 4922
rect 2726 4870 2728 4922
rect 2482 4868 2488 4870
rect 2544 4868 2568 4870
rect 2624 4868 2648 4870
rect 2704 4868 2728 4870
rect 2784 4868 2790 4870
rect 2482 4848 2790 4868
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 2482 3836 2790 3856
rect 2482 3834 2488 3836
rect 2544 3834 2568 3836
rect 2624 3834 2648 3836
rect 2704 3834 2728 3836
rect 2784 3834 2790 3836
rect 2544 3782 2546 3834
rect 2726 3782 2728 3834
rect 2482 3780 2488 3782
rect 2544 3780 2568 3782
rect 2624 3780 2648 3782
rect 2704 3780 2728 3782
rect 2784 3780 2790 3782
rect 2482 3760 2790 3780
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 2240 3482 2268 3538
rect 1780 2990 1808 3470
rect 2240 3454 2360 3482
rect 1846 3292 2154 3312
rect 1846 3290 1852 3292
rect 1908 3290 1932 3292
rect 1988 3290 2012 3292
rect 2068 3290 2092 3292
rect 2148 3290 2154 3292
rect 1908 3238 1910 3290
rect 2090 3238 2092 3290
rect 1846 3236 1852 3238
rect 1908 3236 1932 3238
rect 1988 3236 2012 3238
rect 2068 3236 2092 3238
rect 2148 3236 2154 3238
rect 1846 3216 2154 3236
rect 2332 3194 2360 3454
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 1768 2984 1820 2990
rect 1768 2926 1820 2932
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1688 2514 1716 2790
rect 1676 2508 1728 2514
rect 1676 2450 1728 2456
rect 1676 2372 1728 2378
rect 1676 2314 1728 2320
rect 1688 1426 1716 2314
rect 1780 2310 1808 2926
rect 1860 2848 1912 2854
rect 1860 2790 1912 2796
rect 1872 2378 1900 2790
rect 1860 2372 1912 2378
rect 1860 2314 1912 2320
rect 2228 2372 2280 2378
rect 2228 2314 2280 2320
rect 1768 2304 1820 2310
rect 1768 2246 1820 2252
rect 1676 1420 1728 1426
rect 1676 1362 1728 1368
rect 1780 1222 1808 2246
rect 1846 2204 2154 2224
rect 1846 2202 1852 2204
rect 1908 2202 1932 2204
rect 1988 2202 2012 2204
rect 2068 2202 2092 2204
rect 2148 2202 2154 2204
rect 1908 2150 1910 2202
rect 2090 2150 2092 2202
rect 1846 2148 1852 2150
rect 1908 2148 1932 2150
rect 1988 2148 2012 2150
rect 2068 2148 2092 2150
rect 2148 2148 2154 2150
rect 1846 2128 2154 2148
rect 1860 2032 1912 2038
rect 1860 1974 1912 1980
rect 1872 1562 1900 1974
rect 2044 1896 2096 1902
rect 2044 1838 2096 1844
rect 2056 1562 2084 1838
rect 1860 1556 1912 1562
rect 1860 1498 1912 1504
rect 2044 1556 2096 1562
rect 2044 1498 2096 1504
rect 2240 1494 2268 2314
rect 2332 1970 2360 3130
rect 2482 2748 2790 2768
rect 2482 2746 2488 2748
rect 2544 2746 2568 2748
rect 2624 2746 2648 2748
rect 2704 2746 2728 2748
rect 2784 2746 2790 2748
rect 2544 2694 2546 2746
rect 2726 2694 2728 2746
rect 2482 2692 2488 2694
rect 2544 2692 2568 2694
rect 2624 2692 2648 2694
rect 2704 2692 2728 2694
rect 2784 2692 2790 2694
rect 2482 2672 2790 2692
rect 2412 2644 2464 2650
rect 2412 2586 2464 2592
rect 2320 1964 2372 1970
rect 2320 1906 2372 1912
rect 2228 1488 2280 1494
rect 2228 1430 2280 1436
rect 2424 1290 2452 2586
rect 2884 2038 2912 4014
rect 2976 3602 3004 4626
rect 3514 4448 3570 4457
rect 3118 4380 3426 4400
rect 3514 4383 3570 4392
rect 3118 4378 3124 4380
rect 3180 4378 3204 4380
rect 3260 4378 3284 4380
rect 3340 4378 3364 4380
rect 3420 4378 3426 4380
rect 3180 4326 3182 4378
rect 3362 4326 3364 4378
rect 3118 4324 3124 4326
rect 3180 4324 3204 4326
rect 3260 4324 3284 4326
rect 3340 4324 3364 4326
rect 3420 4324 3426 4326
rect 3118 4304 3426 4324
rect 3528 3942 3556 4383
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 2964 3596 3016 3602
rect 2964 3538 3016 3544
rect 2976 2582 3004 3538
rect 3118 3292 3426 3312
rect 3118 3290 3124 3292
rect 3180 3290 3204 3292
rect 3260 3290 3284 3292
rect 3340 3290 3364 3292
rect 3420 3290 3426 3292
rect 3180 3238 3182 3290
rect 3362 3238 3364 3290
rect 3118 3236 3124 3238
rect 3180 3236 3204 3238
rect 3260 3236 3284 3238
rect 3340 3236 3364 3238
rect 3420 3236 3426 3238
rect 3118 3216 3426 3236
rect 2964 2576 3016 2582
rect 2964 2518 3016 2524
rect 2872 2032 2924 2038
rect 2872 1974 2924 1980
rect 2976 1902 3004 2518
rect 3606 2408 3662 2417
rect 3606 2343 3662 2352
rect 3118 2204 3426 2224
rect 3118 2202 3124 2204
rect 3180 2202 3204 2204
rect 3260 2202 3284 2204
rect 3340 2202 3364 2204
rect 3420 2202 3426 2204
rect 3180 2150 3182 2202
rect 3362 2150 3364 2202
rect 3118 2148 3124 2150
rect 3180 2148 3204 2150
rect 3260 2148 3284 2150
rect 3340 2148 3364 2150
rect 3420 2148 3426 2150
rect 3118 2128 3426 2148
rect 2964 1896 3016 1902
rect 2964 1838 3016 1844
rect 2872 1760 2924 1766
rect 2872 1702 2924 1708
rect 2482 1660 2790 1680
rect 2482 1658 2488 1660
rect 2544 1658 2568 1660
rect 2624 1658 2648 1660
rect 2704 1658 2728 1660
rect 2784 1658 2790 1660
rect 2544 1606 2546 1658
rect 2726 1606 2728 1658
rect 2482 1604 2488 1606
rect 2544 1604 2568 1606
rect 2624 1604 2648 1606
rect 2704 1604 2728 1606
rect 2784 1604 2790 1606
rect 2482 1584 2790 1604
rect 2412 1284 2464 1290
rect 2412 1226 2464 1232
rect 1768 1216 1820 1222
rect 1768 1158 1820 1164
rect 1846 1116 2154 1136
rect 1846 1114 1852 1116
rect 1908 1114 1932 1116
rect 1988 1114 2012 1116
rect 2068 1114 2092 1116
rect 2148 1114 2154 1116
rect 1908 1062 1910 1114
rect 2090 1062 2092 1114
rect 1846 1060 1852 1062
rect 1908 1060 1932 1062
rect 1988 1060 2012 1062
rect 2068 1060 2092 1062
rect 2148 1060 2154 1062
rect 1846 1040 2154 1060
rect 2884 814 2912 1702
rect 3620 1494 3648 2343
rect 3608 1488 3660 1494
rect 3514 1456 3570 1465
rect 3608 1430 3660 1436
rect 3514 1391 3570 1400
rect 3118 1116 3426 1136
rect 3118 1114 3124 1116
rect 3180 1114 3204 1116
rect 3260 1114 3284 1116
rect 3340 1114 3364 1116
rect 3420 1114 3426 1116
rect 3180 1062 3182 1114
rect 3362 1062 3364 1114
rect 3118 1060 3124 1062
rect 3180 1060 3204 1062
rect 3260 1060 3284 1062
rect 3340 1060 3364 1062
rect 3420 1060 3426 1062
rect 3118 1040 3426 1060
rect 3528 1018 3556 1391
rect 3516 1012 3568 1018
rect 3516 954 3568 960
rect 480 808 532 814
rect 480 750 532 756
rect 1584 808 1636 814
rect 1584 750 1636 756
rect 2872 808 2924 814
rect 2872 750 2924 756
rect 2964 740 3016 746
rect 2964 682 3016 688
rect 1210 572 1518 592
rect 1210 570 1216 572
rect 1272 570 1296 572
rect 1352 570 1376 572
rect 1432 570 1456 572
rect 1512 570 1518 572
rect 1272 518 1274 570
rect 1454 518 1456 570
rect 1210 516 1216 518
rect 1272 516 1296 518
rect 1352 516 1376 518
rect 1432 516 1456 518
rect 1512 516 1518 518
rect 1210 496 1518 516
rect 2482 572 2790 592
rect 2482 570 2488 572
rect 2544 570 2568 572
rect 2624 570 2648 572
rect 2704 570 2728 572
rect 2784 570 2790 572
rect 2544 518 2546 570
rect 2726 518 2728 570
rect 2482 516 2488 518
rect 2544 516 2568 518
rect 2624 516 2648 518
rect 2704 516 2728 518
rect 2784 516 2790 518
rect 2482 496 2790 516
rect 2976 513 3004 682
rect 2962 504 3018 513
rect 2962 439 3018 448
<< via2 >>
rect 1950 7184 2006 7240
rect 1216 7098 1272 7100
rect 1296 7098 1352 7100
rect 1376 7098 1432 7100
rect 1456 7098 1512 7100
rect 1216 7046 1262 7098
rect 1262 7046 1272 7098
rect 1296 7046 1326 7098
rect 1326 7046 1338 7098
rect 1338 7046 1352 7098
rect 1376 7046 1390 7098
rect 1390 7046 1402 7098
rect 1402 7046 1432 7098
rect 1456 7046 1466 7098
rect 1466 7046 1512 7098
rect 1216 7044 1272 7046
rect 1296 7044 1352 7046
rect 1376 7044 1432 7046
rect 1456 7044 1512 7046
rect 2488 7098 2544 7100
rect 2568 7098 2624 7100
rect 2648 7098 2704 7100
rect 2728 7098 2784 7100
rect 2488 7046 2534 7098
rect 2534 7046 2544 7098
rect 2568 7046 2598 7098
rect 2598 7046 2610 7098
rect 2610 7046 2624 7098
rect 2648 7046 2662 7098
rect 2662 7046 2674 7098
rect 2674 7046 2704 7098
rect 2728 7046 2738 7098
rect 2738 7046 2784 7098
rect 2488 7044 2544 7046
rect 2568 7044 2624 7046
rect 2648 7044 2704 7046
rect 2728 7044 2784 7046
rect 294 6568 350 6624
rect 580 6554 636 6556
rect 660 6554 716 6556
rect 740 6554 796 6556
rect 820 6554 876 6556
rect 580 6502 626 6554
rect 626 6502 636 6554
rect 660 6502 690 6554
rect 690 6502 702 6554
rect 702 6502 716 6554
rect 740 6502 754 6554
rect 754 6502 766 6554
rect 766 6502 796 6554
rect 820 6502 830 6554
rect 830 6502 876 6554
rect 580 6500 636 6502
rect 660 6500 716 6502
rect 740 6500 796 6502
rect 820 6500 876 6502
rect 1852 6554 1908 6556
rect 1932 6554 1988 6556
rect 2012 6554 2068 6556
rect 2092 6554 2148 6556
rect 1852 6502 1898 6554
rect 1898 6502 1908 6554
rect 1932 6502 1962 6554
rect 1962 6502 1974 6554
rect 1974 6502 1988 6554
rect 2012 6502 2026 6554
rect 2026 6502 2038 6554
rect 2038 6502 2068 6554
rect 2092 6502 2102 6554
rect 2102 6502 2148 6554
rect 1852 6500 1908 6502
rect 1932 6500 1988 6502
rect 2012 6500 2068 6502
rect 2092 6500 2148 6502
rect 1216 6010 1272 6012
rect 1296 6010 1352 6012
rect 1376 6010 1432 6012
rect 1456 6010 1512 6012
rect 1216 5958 1262 6010
rect 1262 5958 1272 6010
rect 1296 5958 1326 6010
rect 1326 5958 1338 6010
rect 1338 5958 1352 6010
rect 1376 5958 1390 6010
rect 1390 5958 1402 6010
rect 1402 5958 1432 6010
rect 1456 5958 1466 6010
rect 1466 5958 1512 6010
rect 1216 5956 1272 5958
rect 1296 5956 1352 5958
rect 1376 5956 1432 5958
rect 1456 5956 1512 5958
rect 580 5466 636 5468
rect 660 5466 716 5468
rect 740 5466 796 5468
rect 820 5466 876 5468
rect 580 5414 626 5466
rect 626 5414 636 5466
rect 660 5414 690 5466
rect 690 5414 702 5466
rect 702 5414 716 5466
rect 740 5414 754 5466
rect 754 5414 766 5466
rect 766 5414 796 5466
rect 820 5414 830 5466
rect 830 5414 876 5466
rect 580 5412 636 5414
rect 660 5412 716 5414
rect 740 5412 796 5414
rect 820 5412 876 5414
rect 580 4378 636 4380
rect 660 4378 716 4380
rect 740 4378 796 4380
rect 820 4378 876 4380
rect 580 4326 626 4378
rect 626 4326 636 4378
rect 660 4326 690 4378
rect 690 4326 702 4378
rect 702 4326 716 4378
rect 740 4326 754 4378
rect 754 4326 766 4378
rect 766 4326 796 4378
rect 820 4326 830 4378
rect 830 4326 876 4378
rect 580 4324 636 4326
rect 660 4324 716 4326
rect 740 4324 796 4326
rect 820 4324 876 4326
rect 478 3848 534 3904
rect 580 3290 636 3292
rect 660 3290 716 3292
rect 740 3290 796 3292
rect 820 3290 876 3292
rect 580 3238 626 3290
rect 626 3238 636 3290
rect 660 3238 690 3290
rect 690 3238 702 3290
rect 702 3238 716 3290
rect 740 3238 754 3290
rect 754 3238 766 3290
rect 766 3238 796 3290
rect 820 3238 830 3290
rect 830 3238 876 3290
rect 580 3236 636 3238
rect 660 3236 716 3238
rect 740 3236 796 3238
rect 820 3236 876 3238
rect 1216 4922 1272 4924
rect 1296 4922 1352 4924
rect 1376 4922 1432 4924
rect 1456 4922 1512 4924
rect 1216 4870 1262 4922
rect 1262 4870 1272 4922
rect 1296 4870 1326 4922
rect 1326 4870 1338 4922
rect 1338 4870 1352 4922
rect 1376 4870 1390 4922
rect 1390 4870 1402 4922
rect 1402 4870 1432 4922
rect 1456 4870 1466 4922
rect 1466 4870 1512 4922
rect 1216 4868 1272 4870
rect 1296 4868 1352 4870
rect 1376 4868 1432 4870
rect 1456 4868 1512 4870
rect 1216 3834 1272 3836
rect 1296 3834 1352 3836
rect 1376 3834 1432 3836
rect 1456 3834 1512 3836
rect 1216 3782 1262 3834
rect 1262 3782 1272 3834
rect 1296 3782 1326 3834
rect 1326 3782 1338 3834
rect 1338 3782 1352 3834
rect 1376 3782 1390 3834
rect 1390 3782 1402 3834
rect 1402 3782 1432 3834
rect 1456 3782 1466 3834
rect 1466 3782 1512 3834
rect 1216 3780 1272 3782
rect 1296 3780 1352 3782
rect 1376 3780 1432 3782
rect 1456 3780 1512 3782
rect 580 2202 636 2204
rect 660 2202 716 2204
rect 740 2202 796 2204
rect 820 2202 876 2204
rect 580 2150 626 2202
rect 626 2150 636 2202
rect 660 2150 690 2202
rect 690 2150 702 2202
rect 702 2150 716 2202
rect 740 2150 754 2202
rect 754 2150 766 2202
rect 766 2150 796 2202
rect 820 2150 830 2202
rect 830 2150 876 2202
rect 580 2148 636 2150
rect 660 2148 716 2150
rect 740 2148 796 2150
rect 820 2148 876 2150
rect 1398 3440 1454 3496
rect 1216 2746 1272 2748
rect 1296 2746 1352 2748
rect 1376 2746 1432 2748
rect 1456 2746 1512 2748
rect 1216 2694 1262 2746
rect 1262 2694 1272 2746
rect 1296 2694 1326 2746
rect 1326 2694 1338 2746
rect 1338 2694 1352 2746
rect 1376 2694 1390 2746
rect 1390 2694 1402 2746
rect 1402 2694 1432 2746
rect 1456 2694 1466 2746
rect 1466 2694 1512 2746
rect 1216 2692 1272 2694
rect 1296 2692 1352 2694
rect 1376 2692 1432 2694
rect 1456 2692 1512 2694
rect 1216 1658 1272 1660
rect 1296 1658 1352 1660
rect 1376 1658 1432 1660
rect 1456 1658 1512 1660
rect 1216 1606 1262 1658
rect 1262 1606 1272 1658
rect 1296 1606 1326 1658
rect 1326 1606 1338 1658
rect 1338 1606 1352 1658
rect 1376 1606 1390 1658
rect 1390 1606 1402 1658
rect 1402 1606 1432 1658
rect 1456 1606 1466 1658
rect 1466 1606 1512 1658
rect 1216 1604 1272 1606
rect 1296 1604 1352 1606
rect 1376 1604 1432 1606
rect 1456 1604 1512 1606
rect 478 1264 534 1320
rect 580 1114 636 1116
rect 660 1114 716 1116
rect 740 1114 796 1116
rect 820 1114 876 1116
rect 580 1062 626 1114
rect 626 1062 636 1114
rect 660 1062 690 1114
rect 690 1062 702 1114
rect 702 1062 716 1114
rect 740 1062 754 1114
rect 754 1062 766 1114
rect 766 1062 796 1114
rect 820 1062 830 1114
rect 830 1062 876 1114
rect 580 1060 636 1062
rect 660 1060 716 1062
rect 740 1060 796 1062
rect 820 1060 876 1062
rect 1852 5466 1908 5468
rect 1932 5466 1988 5468
rect 2012 5466 2068 5468
rect 2092 5466 2148 5468
rect 1852 5414 1898 5466
rect 1898 5414 1908 5466
rect 1932 5414 1962 5466
rect 1962 5414 1974 5466
rect 1974 5414 1988 5466
rect 2012 5414 2026 5466
rect 2026 5414 2038 5466
rect 2038 5414 2068 5466
rect 2092 5414 2102 5466
rect 2102 5414 2148 5466
rect 1852 5412 1908 5414
rect 1932 5412 1988 5414
rect 2012 5412 2068 5414
rect 2092 5412 2148 5414
rect 3124 6554 3180 6556
rect 3204 6554 3260 6556
rect 3284 6554 3340 6556
rect 3364 6554 3420 6556
rect 3124 6502 3170 6554
rect 3170 6502 3180 6554
rect 3204 6502 3234 6554
rect 3234 6502 3246 6554
rect 3246 6502 3260 6554
rect 3284 6502 3298 6554
rect 3298 6502 3310 6554
rect 3310 6502 3340 6554
rect 3364 6502 3374 6554
rect 3374 6502 3420 6554
rect 3124 6500 3180 6502
rect 3204 6500 3260 6502
rect 3284 6500 3340 6502
rect 3364 6500 3420 6502
rect 3514 6432 3570 6488
rect 1852 4378 1908 4380
rect 1932 4378 1988 4380
rect 2012 4378 2068 4380
rect 2092 4378 2148 4380
rect 1852 4326 1898 4378
rect 1898 4326 1908 4378
rect 1932 4326 1962 4378
rect 1962 4326 1974 4378
rect 1974 4326 1988 4378
rect 2012 4326 2026 4378
rect 2026 4326 2038 4378
rect 2038 4326 2068 4378
rect 2092 4326 2102 4378
rect 2102 4326 2148 4378
rect 1852 4324 1908 4326
rect 1932 4324 1988 4326
rect 2012 4324 2068 4326
rect 2092 4324 2148 4326
rect 2488 6010 2544 6012
rect 2568 6010 2624 6012
rect 2648 6010 2704 6012
rect 2728 6010 2784 6012
rect 2488 5958 2534 6010
rect 2534 5958 2544 6010
rect 2568 5958 2598 6010
rect 2598 5958 2610 6010
rect 2610 5958 2624 6010
rect 2648 5958 2662 6010
rect 2662 5958 2674 6010
rect 2674 5958 2704 6010
rect 2728 5958 2738 6010
rect 2738 5958 2784 6010
rect 2488 5956 2544 5958
rect 2568 5956 2624 5958
rect 2648 5956 2704 5958
rect 2728 5956 2784 5958
rect 3124 5466 3180 5468
rect 3204 5466 3260 5468
rect 3284 5466 3340 5468
rect 3364 5466 3420 5468
rect 3124 5414 3170 5466
rect 3170 5414 3180 5466
rect 3204 5414 3234 5466
rect 3234 5414 3246 5466
rect 3246 5414 3260 5466
rect 3284 5414 3298 5466
rect 3298 5414 3310 5466
rect 3310 5414 3340 5466
rect 3364 5414 3374 5466
rect 3374 5414 3420 5466
rect 3124 5412 3180 5414
rect 3204 5412 3260 5414
rect 3284 5412 3340 5414
rect 3364 5412 3420 5414
rect 3514 5344 3570 5400
rect 2488 4922 2544 4924
rect 2568 4922 2624 4924
rect 2648 4922 2704 4924
rect 2728 4922 2784 4924
rect 2488 4870 2534 4922
rect 2534 4870 2544 4922
rect 2568 4870 2598 4922
rect 2598 4870 2610 4922
rect 2610 4870 2624 4922
rect 2648 4870 2662 4922
rect 2662 4870 2674 4922
rect 2674 4870 2704 4922
rect 2728 4870 2738 4922
rect 2738 4870 2784 4922
rect 2488 4868 2544 4870
rect 2568 4868 2624 4870
rect 2648 4868 2704 4870
rect 2728 4868 2784 4870
rect 2488 3834 2544 3836
rect 2568 3834 2624 3836
rect 2648 3834 2704 3836
rect 2728 3834 2784 3836
rect 2488 3782 2534 3834
rect 2534 3782 2544 3834
rect 2568 3782 2598 3834
rect 2598 3782 2610 3834
rect 2610 3782 2624 3834
rect 2648 3782 2662 3834
rect 2662 3782 2674 3834
rect 2674 3782 2704 3834
rect 2728 3782 2738 3834
rect 2738 3782 2784 3834
rect 2488 3780 2544 3782
rect 2568 3780 2624 3782
rect 2648 3780 2704 3782
rect 2728 3780 2784 3782
rect 1852 3290 1908 3292
rect 1932 3290 1988 3292
rect 2012 3290 2068 3292
rect 2092 3290 2148 3292
rect 1852 3238 1898 3290
rect 1898 3238 1908 3290
rect 1932 3238 1962 3290
rect 1962 3238 1974 3290
rect 1974 3238 1988 3290
rect 2012 3238 2026 3290
rect 2026 3238 2038 3290
rect 2038 3238 2068 3290
rect 2092 3238 2102 3290
rect 2102 3238 2148 3290
rect 1852 3236 1908 3238
rect 1932 3236 1988 3238
rect 2012 3236 2068 3238
rect 2092 3236 2148 3238
rect 1852 2202 1908 2204
rect 1932 2202 1988 2204
rect 2012 2202 2068 2204
rect 2092 2202 2148 2204
rect 1852 2150 1898 2202
rect 1898 2150 1908 2202
rect 1932 2150 1962 2202
rect 1962 2150 1974 2202
rect 1974 2150 1988 2202
rect 2012 2150 2026 2202
rect 2026 2150 2038 2202
rect 2038 2150 2068 2202
rect 2092 2150 2102 2202
rect 2102 2150 2148 2202
rect 1852 2148 1908 2150
rect 1932 2148 1988 2150
rect 2012 2148 2068 2150
rect 2092 2148 2148 2150
rect 2488 2746 2544 2748
rect 2568 2746 2624 2748
rect 2648 2746 2704 2748
rect 2728 2746 2784 2748
rect 2488 2694 2534 2746
rect 2534 2694 2544 2746
rect 2568 2694 2598 2746
rect 2598 2694 2610 2746
rect 2610 2694 2624 2746
rect 2648 2694 2662 2746
rect 2662 2694 2674 2746
rect 2674 2694 2704 2746
rect 2728 2694 2738 2746
rect 2738 2694 2784 2746
rect 2488 2692 2544 2694
rect 2568 2692 2624 2694
rect 2648 2692 2704 2694
rect 2728 2692 2784 2694
rect 3514 4392 3570 4448
rect 3124 4378 3180 4380
rect 3204 4378 3260 4380
rect 3284 4378 3340 4380
rect 3364 4378 3420 4380
rect 3124 4326 3170 4378
rect 3170 4326 3180 4378
rect 3204 4326 3234 4378
rect 3234 4326 3246 4378
rect 3246 4326 3260 4378
rect 3284 4326 3298 4378
rect 3298 4326 3310 4378
rect 3310 4326 3340 4378
rect 3364 4326 3374 4378
rect 3374 4326 3420 4378
rect 3124 4324 3180 4326
rect 3204 4324 3260 4326
rect 3284 4324 3340 4326
rect 3364 4324 3420 4326
rect 3124 3290 3180 3292
rect 3204 3290 3260 3292
rect 3284 3290 3340 3292
rect 3364 3290 3420 3292
rect 3124 3238 3170 3290
rect 3170 3238 3180 3290
rect 3204 3238 3234 3290
rect 3234 3238 3246 3290
rect 3246 3238 3260 3290
rect 3284 3238 3298 3290
rect 3298 3238 3310 3290
rect 3310 3238 3340 3290
rect 3364 3238 3374 3290
rect 3374 3238 3420 3290
rect 3124 3236 3180 3238
rect 3204 3236 3260 3238
rect 3284 3236 3340 3238
rect 3364 3236 3420 3238
rect 3606 2352 3662 2408
rect 3124 2202 3180 2204
rect 3204 2202 3260 2204
rect 3284 2202 3340 2204
rect 3364 2202 3420 2204
rect 3124 2150 3170 2202
rect 3170 2150 3180 2202
rect 3204 2150 3234 2202
rect 3234 2150 3246 2202
rect 3246 2150 3260 2202
rect 3284 2150 3298 2202
rect 3298 2150 3310 2202
rect 3310 2150 3340 2202
rect 3364 2150 3374 2202
rect 3374 2150 3420 2202
rect 3124 2148 3180 2150
rect 3204 2148 3260 2150
rect 3284 2148 3340 2150
rect 3364 2148 3420 2150
rect 2488 1658 2544 1660
rect 2568 1658 2624 1660
rect 2648 1658 2704 1660
rect 2728 1658 2784 1660
rect 2488 1606 2534 1658
rect 2534 1606 2544 1658
rect 2568 1606 2598 1658
rect 2598 1606 2610 1658
rect 2610 1606 2624 1658
rect 2648 1606 2662 1658
rect 2662 1606 2674 1658
rect 2674 1606 2704 1658
rect 2728 1606 2738 1658
rect 2738 1606 2784 1658
rect 2488 1604 2544 1606
rect 2568 1604 2624 1606
rect 2648 1604 2704 1606
rect 2728 1604 2784 1606
rect 1852 1114 1908 1116
rect 1932 1114 1988 1116
rect 2012 1114 2068 1116
rect 2092 1114 2148 1116
rect 1852 1062 1898 1114
rect 1898 1062 1908 1114
rect 1932 1062 1962 1114
rect 1962 1062 1974 1114
rect 1974 1062 1988 1114
rect 2012 1062 2026 1114
rect 2026 1062 2038 1114
rect 2038 1062 2068 1114
rect 2092 1062 2102 1114
rect 2102 1062 2148 1114
rect 1852 1060 1908 1062
rect 1932 1060 1988 1062
rect 2012 1060 2068 1062
rect 2092 1060 2148 1062
rect 3514 1400 3570 1456
rect 3124 1114 3180 1116
rect 3204 1114 3260 1116
rect 3284 1114 3340 1116
rect 3364 1114 3420 1116
rect 3124 1062 3170 1114
rect 3170 1062 3180 1114
rect 3204 1062 3234 1114
rect 3234 1062 3246 1114
rect 3246 1062 3260 1114
rect 3284 1062 3298 1114
rect 3298 1062 3310 1114
rect 3310 1062 3340 1114
rect 3364 1062 3374 1114
rect 3374 1062 3420 1114
rect 3124 1060 3180 1062
rect 3204 1060 3260 1062
rect 3284 1060 3340 1062
rect 3364 1060 3420 1062
rect 1216 570 1272 572
rect 1296 570 1352 572
rect 1376 570 1432 572
rect 1456 570 1512 572
rect 1216 518 1262 570
rect 1262 518 1272 570
rect 1296 518 1326 570
rect 1326 518 1338 570
rect 1338 518 1352 570
rect 1376 518 1390 570
rect 1390 518 1402 570
rect 1402 518 1432 570
rect 1456 518 1466 570
rect 1466 518 1512 570
rect 1216 516 1272 518
rect 1296 516 1352 518
rect 1376 516 1432 518
rect 1456 516 1512 518
rect 2488 570 2544 572
rect 2568 570 2624 572
rect 2648 570 2704 572
rect 2728 570 2784 572
rect 2488 518 2534 570
rect 2534 518 2544 570
rect 2568 518 2598 570
rect 2598 518 2610 570
rect 2610 518 2624 570
rect 2648 518 2662 570
rect 2662 518 2674 570
rect 2674 518 2704 570
rect 2728 518 2738 570
rect 2738 518 2784 570
rect 2488 516 2544 518
rect 2568 516 2624 518
rect 2648 516 2704 518
rect 2728 516 2784 518
rect 2962 448 3018 504
<< metal3 >>
rect 1945 7242 2011 7245
rect 1945 7240 4000 7242
rect 1945 7184 1950 7240
rect 2006 7184 4000 7240
rect 1945 7182 4000 7184
rect 1945 7179 2011 7182
rect 1204 7104 1524 7105
rect 1204 7040 1212 7104
rect 1276 7040 1292 7104
rect 1356 7040 1372 7104
rect 1436 7040 1452 7104
rect 1516 7040 1524 7104
rect 1204 7039 1524 7040
rect 2476 7104 2796 7105
rect 2476 7040 2484 7104
rect 2548 7040 2564 7104
rect 2628 7040 2644 7104
rect 2708 7040 2724 7104
rect 2788 7040 2796 7104
rect 2476 7039 2796 7040
rect 289 6626 355 6629
rect 0 6624 355 6626
rect 0 6568 294 6624
rect 350 6568 355 6624
rect 0 6566 355 6568
rect 289 6563 355 6566
rect 568 6560 888 6561
rect 568 6496 576 6560
rect 640 6496 656 6560
rect 720 6496 736 6560
rect 800 6496 816 6560
rect 880 6496 888 6560
rect 568 6495 888 6496
rect 1840 6560 2160 6561
rect 1840 6496 1848 6560
rect 1912 6496 1928 6560
rect 1992 6496 2008 6560
rect 2072 6496 2088 6560
rect 2152 6496 2160 6560
rect 1840 6495 2160 6496
rect 3112 6560 3432 6561
rect 3112 6496 3120 6560
rect 3184 6496 3200 6560
rect 3264 6496 3280 6560
rect 3344 6496 3360 6560
rect 3424 6496 3432 6560
rect 3112 6495 3432 6496
rect 3509 6490 3575 6493
rect 3509 6488 4000 6490
rect 3509 6432 3514 6488
rect 3570 6432 4000 6488
rect 3509 6430 4000 6432
rect 3509 6427 3575 6430
rect 1204 6016 1524 6017
rect 1204 5952 1212 6016
rect 1276 5952 1292 6016
rect 1356 5952 1372 6016
rect 1436 5952 1452 6016
rect 1516 5952 1524 6016
rect 1204 5951 1524 5952
rect 2476 6016 2796 6017
rect 2476 5952 2484 6016
rect 2548 5952 2564 6016
rect 2628 5952 2644 6016
rect 2708 5952 2724 6016
rect 2788 5952 2796 6016
rect 2476 5951 2796 5952
rect 568 5472 888 5473
rect 568 5408 576 5472
rect 640 5408 656 5472
rect 720 5408 736 5472
rect 800 5408 816 5472
rect 880 5408 888 5472
rect 568 5407 888 5408
rect 1840 5472 2160 5473
rect 1840 5408 1848 5472
rect 1912 5408 1928 5472
rect 1992 5408 2008 5472
rect 2072 5408 2088 5472
rect 2152 5408 2160 5472
rect 1840 5407 2160 5408
rect 3112 5472 3432 5473
rect 3112 5408 3120 5472
rect 3184 5408 3200 5472
rect 3264 5408 3280 5472
rect 3344 5408 3360 5472
rect 3424 5408 3432 5472
rect 3112 5407 3432 5408
rect 3509 5402 3575 5405
rect 3509 5400 4000 5402
rect 3509 5344 3514 5400
rect 3570 5344 4000 5400
rect 3509 5342 4000 5344
rect 3509 5339 3575 5342
rect 1204 4928 1524 4929
rect 1204 4864 1212 4928
rect 1276 4864 1292 4928
rect 1356 4864 1372 4928
rect 1436 4864 1452 4928
rect 1516 4864 1524 4928
rect 1204 4863 1524 4864
rect 2476 4928 2796 4929
rect 2476 4864 2484 4928
rect 2548 4864 2564 4928
rect 2628 4864 2644 4928
rect 2708 4864 2724 4928
rect 2788 4864 2796 4928
rect 2476 4863 2796 4864
rect 3509 4450 3575 4453
rect 3509 4448 4000 4450
rect 3509 4392 3514 4448
rect 3570 4392 4000 4448
rect 3509 4390 4000 4392
rect 3509 4387 3575 4390
rect 568 4384 888 4385
rect 568 4320 576 4384
rect 640 4320 656 4384
rect 720 4320 736 4384
rect 800 4320 816 4384
rect 880 4320 888 4384
rect 568 4319 888 4320
rect 1840 4384 2160 4385
rect 1840 4320 1848 4384
rect 1912 4320 1928 4384
rect 1992 4320 2008 4384
rect 2072 4320 2088 4384
rect 2152 4320 2160 4384
rect 1840 4319 2160 4320
rect 3112 4384 3432 4385
rect 3112 4320 3120 4384
rect 3184 4320 3200 4384
rect 3264 4320 3280 4384
rect 3344 4320 3360 4384
rect 3424 4320 3432 4384
rect 3112 4319 3432 4320
rect 473 3906 539 3909
rect 0 3904 539 3906
rect 0 3848 478 3904
rect 534 3848 539 3904
rect 0 3846 539 3848
rect 473 3843 539 3846
rect 1204 3840 1524 3841
rect 1204 3776 1212 3840
rect 1276 3776 1292 3840
rect 1356 3776 1372 3840
rect 1436 3776 1452 3840
rect 1516 3776 1524 3840
rect 1204 3775 1524 3776
rect 2476 3840 2796 3841
rect 2476 3776 2484 3840
rect 2548 3776 2564 3840
rect 2628 3776 2644 3840
rect 2708 3776 2724 3840
rect 2788 3776 2796 3840
rect 2476 3775 2796 3776
rect 1393 3498 1459 3501
rect 1393 3496 4000 3498
rect 1393 3440 1398 3496
rect 1454 3440 4000 3496
rect 1393 3438 4000 3440
rect 1393 3435 1459 3438
rect 568 3296 888 3297
rect 568 3232 576 3296
rect 640 3232 656 3296
rect 720 3232 736 3296
rect 800 3232 816 3296
rect 880 3232 888 3296
rect 568 3231 888 3232
rect 1840 3296 2160 3297
rect 1840 3232 1848 3296
rect 1912 3232 1928 3296
rect 1992 3232 2008 3296
rect 2072 3232 2088 3296
rect 2152 3232 2160 3296
rect 1840 3231 2160 3232
rect 3112 3296 3432 3297
rect 3112 3232 3120 3296
rect 3184 3232 3200 3296
rect 3264 3232 3280 3296
rect 3344 3232 3360 3296
rect 3424 3232 3432 3296
rect 3112 3231 3432 3232
rect 1204 2752 1524 2753
rect 1204 2688 1212 2752
rect 1276 2688 1292 2752
rect 1356 2688 1372 2752
rect 1436 2688 1452 2752
rect 1516 2688 1524 2752
rect 1204 2687 1524 2688
rect 2476 2752 2796 2753
rect 2476 2688 2484 2752
rect 2548 2688 2564 2752
rect 2628 2688 2644 2752
rect 2708 2688 2724 2752
rect 2788 2688 2796 2752
rect 2476 2687 2796 2688
rect 3601 2410 3667 2413
rect 3601 2408 4000 2410
rect 3601 2352 3606 2408
rect 3662 2352 4000 2408
rect 3601 2350 4000 2352
rect 3601 2347 3667 2350
rect 568 2208 888 2209
rect 568 2144 576 2208
rect 640 2144 656 2208
rect 720 2144 736 2208
rect 800 2144 816 2208
rect 880 2144 888 2208
rect 568 2143 888 2144
rect 1840 2208 2160 2209
rect 1840 2144 1848 2208
rect 1912 2144 1928 2208
rect 1992 2144 2008 2208
rect 2072 2144 2088 2208
rect 2152 2144 2160 2208
rect 1840 2143 2160 2144
rect 3112 2208 3432 2209
rect 3112 2144 3120 2208
rect 3184 2144 3200 2208
rect 3264 2144 3280 2208
rect 3344 2144 3360 2208
rect 3424 2144 3432 2208
rect 3112 2143 3432 2144
rect 1204 1664 1524 1665
rect 1204 1600 1212 1664
rect 1276 1600 1292 1664
rect 1356 1600 1372 1664
rect 1436 1600 1452 1664
rect 1516 1600 1524 1664
rect 1204 1599 1524 1600
rect 2476 1664 2796 1665
rect 2476 1600 2484 1664
rect 2548 1600 2564 1664
rect 2628 1600 2644 1664
rect 2708 1600 2724 1664
rect 2788 1600 2796 1664
rect 2476 1599 2796 1600
rect 3509 1458 3575 1461
rect 3509 1456 4000 1458
rect 3509 1400 3514 1456
rect 3570 1400 4000 1456
rect 3509 1398 4000 1400
rect 3509 1395 3575 1398
rect 473 1322 539 1325
rect 0 1320 539 1322
rect 0 1264 478 1320
rect 534 1264 539 1320
rect 0 1262 539 1264
rect 473 1259 539 1262
rect 568 1120 888 1121
rect 568 1056 576 1120
rect 640 1056 656 1120
rect 720 1056 736 1120
rect 800 1056 816 1120
rect 880 1056 888 1120
rect 568 1055 888 1056
rect 1840 1120 2160 1121
rect 1840 1056 1848 1120
rect 1912 1056 1928 1120
rect 1992 1056 2008 1120
rect 2072 1056 2088 1120
rect 2152 1056 2160 1120
rect 1840 1055 2160 1056
rect 3112 1120 3432 1121
rect 3112 1056 3120 1120
rect 3184 1056 3200 1120
rect 3264 1056 3280 1120
rect 3344 1056 3360 1120
rect 3424 1056 3432 1120
rect 3112 1055 3432 1056
rect 1204 576 1524 577
rect 1204 512 1212 576
rect 1276 512 1292 576
rect 1356 512 1372 576
rect 1436 512 1452 576
rect 1516 512 1524 576
rect 1204 511 1524 512
rect 2476 576 2796 577
rect 2476 512 2484 576
rect 2548 512 2564 576
rect 2628 512 2644 576
rect 2708 512 2724 576
rect 2788 512 2796 576
rect 2476 511 2796 512
rect 2957 506 3023 509
rect 2957 504 4000 506
rect 2957 448 2962 504
rect 3018 448 4000 504
rect 2957 446 4000 448
rect 2957 443 3023 446
<< via3 >>
rect 1212 7100 1276 7104
rect 1212 7044 1216 7100
rect 1216 7044 1272 7100
rect 1272 7044 1276 7100
rect 1212 7040 1276 7044
rect 1292 7100 1356 7104
rect 1292 7044 1296 7100
rect 1296 7044 1352 7100
rect 1352 7044 1356 7100
rect 1292 7040 1356 7044
rect 1372 7100 1436 7104
rect 1372 7044 1376 7100
rect 1376 7044 1432 7100
rect 1432 7044 1436 7100
rect 1372 7040 1436 7044
rect 1452 7100 1516 7104
rect 1452 7044 1456 7100
rect 1456 7044 1512 7100
rect 1512 7044 1516 7100
rect 1452 7040 1516 7044
rect 2484 7100 2548 7104
rect 2484 7044 2488 7100
rect 2488 7044 2544 7100
rect 2544 7044 2548 7100
rect 2484 7040 2548 7044
rect 2564 7100 2628 7104
rect 2564 7044 2568 7100
rect 2568 7044 2624 7100
rect 2624 7044 2628 7100
rect 2564 7040 2628 7044
rect 2644 7100 2708 7104
rect 2644 7044 2648 7100
rect 2648 7044 2704 7100
rect 2704 7044 2708 7100
rect 2644 7040 2708 7044
rect 2724 7100 2788 7104
rect 2724 7044 2728 7100
rect 2728 7044 2784 7100
rect 2784 7044 2788 7100
rect 2724 7040 2788 7044
rect 576 6556 640 6560
rect 576 6500 580 6556
rect 580 6500 636 6556
rect 636 6500 640 6556
rect 576 6496 640 6500
rect 656 6556 720 6560
rect 656 6500 660 6556
rect 660 6500 716 6556
rect 716 6500 720 6556
rect 656 6496 720 6500
rect 736 6556 800 6560
rect 736 6500 740 6556
rect 740 6500 796 6556
rect 796 6500 800 6556
rect 736 6496 800 6500
rect 816 6556 880 6560
rect 816 6500 820 6556
rect 820 6500 876 6556
rect 876 6500 880 6556
rect 816 6496 880 6500
rect 1848 6556 1912 6560
rect 1848 6500 1852 6556
rect 1852 6500 1908 6556
rect 1908 6500 1912 6556
rect 1848 6496 1912 6500
rect 1928 6556 1992 6560
rect 1928 6500 1932 6556
rect 1932 6500 1988 6556
rect 1988 6500 1992 6556
rect 1928 6496 1992 6500
rect 2008 6556 2072 6560
rect 2008 6500 2012 6556
rect 2012 6500 2068 6556
rect 2068 6500 2072 6556
rect 2008 6496 2072 6500
rect 2088 6556 2152 6560
rect 2088 6500 2092 6556
rect 2092 6500 2148 6556
rect 2148 6500 2152 6556
rect 2088 6496 2152 6500
rect 3120 6556 3184 6560
rect 3120 6500 3124 6556
rect 3124 6500 3180 6556
rect 3180 6500 3184 6556
rect 3120 6496 3184 6500
rect 3200 6556 3264 6560
rect 3200 6500 3204 6556
rect 3204 6500 3260 6556
rect 3260 6500 3264 6556
rect 3200 6496 3264 6500
rect 3280 6556 3344 6560
rect 3280 6500 3284 6556
rect 3284 6500 3340 6556
rect 3340 6500 3344 6556
rect 3280 6496 3344 6500
rect 3360 6556 3424 6560
rect 3360 6500 3364 6556
rect 3364 6500 3420 6556
rect 3420 6500 3424 6556
rect 3360 6496 3424 6500
rect 1212 6012 1276 6016
rect 1212 5956 1216 6012
rect 1216 5956 1272 6012
rect 1272 5956 1276 6012
rect 1212 5952 1276 5956
rect 1292 6012 1356 6016
rect 1292 5956 1296 6012
rect 1296 5956 1352 6012
rect 1352 5956 1356 6012
rect 1292 5952 1356 5956
rect 1372 6012 1436 6016
rect 1372 5956 1376 6012
rect 1376 5956 1432 6012
rect 1432 5956 1436 6012
rect 1372 5952 1436 5956
rect 1452 6012 1516 6016
rect 1452 5956 1456 6012
rect 1456 5956 1512 6012
rect 1512 5956 1516 6012
rect 1452 5952 1516 5956
rect 2484 6012 2548 6016
rect 2484 5956 2488 6012
rect 2488 5956 2544 6012
rect 2544 5956 2548 6012
rect 2484 5952 2548 5956
rect 2564 6012 2628 6016
rect 2564 5956 2568 6012
rect 2568 5956 2624 6012
rect 2624 5956 2628 6012
rect 2564 5952 2628 5956
rect 2644 6012 2708 6016
rect 2644 5956 2648 6012
rect 2648 5956 2704 6012
rect 2704 5956 2708 6012
rect 2644 5952 2708 5956
rect 2724 6012 2788 6016
rect 2724 5956 2728 6012
rect 2728 5956 2784 6012
rect 2784 5956 2788 6012
rect 2724 5952 2788 5956
rect 576 5468 640 5472
rect 576 5412 580 5468
rect 580 5412 636 5468
rect 636 5412 640 5468
rect 576 5408 640 5412
rect 656 5468 720 5472
rect 656 5412 660 5468
rect 660 5412 716 5468
rect 716 5412 720 5468
rect 656 5408 720 5412
rect 736 5468 800 5472
rect 736 5412 740 5468
rect 740 5412 796 5468
rect 796 5412 800 5468
rect 736 5408 800 5412
rect 816 5468 880 5472
rect 816 5412 820 5468
rect 820 5412 876 5468
rect 876 5412 880 5468
rect 816 5408 880 5412
rect 1848 5468 1912 5472
rect 1848 5412 1852 5468
rect 1852 5412 1908 5468
rect 1908 5412 1912 5468
rect 1848 5408 1912 5412
rect 1928 5468 1992 5472
rect 1928 5412 1932 5468
rect 1932 5412 1988 5468
rect 1988 5412 1992 5468
rect 1928 5408 1992 5412
rect 2008 5468 2072 5472
rect 2008 5412 2012 5468
rect 2012 5412 2068 5468
rect 2068 5412 2072 5468
rect 2008 5408 2072 5412
rect 2088 5468 2152 5472
rect 2088 5412 2092 5468
rect 2092 5412 2148 5468
rect 2148 5412 2152 5468
rect 2088 5408 2152 5412
rect 3120 5468 3184 5472
rect 3120 5412 3124 5468
rect 3124 5412 3180 5468
rect 3180 5412 3184 5468
rect 3120 5408 3184 5412
rect 3200 5468 3264 5472
rect 3200 5412 3204 5468
rect 3204 5412 3260 5468
rect 3260 5412 3264 5468
rect 3200 5408 3264 5412
rect 3280 5468 3344 5472
rect 3280 5412 3284 5468
rect 3284 5412 3340 5468
rect 3340 5412 3344 5468
rect 3280 5408 3344 5412
rect 3360 5468 3424 5472
rect 3360 5412 3364 5468
rect 3364 5412 3420 5468
rect 3420 5412 3424 5468
rect 3360 5408 3424 5412
rect 1212 4924 1276 4928
rect 1212 4868 1216 4924
rect 1216 4868 1272 4924
rect 1272 4868 1276 4924
rect 1212 4864 1276 4868
rect 1292 4924 1356 4928
rect 1292 4868 1296 4924
rect 1296 4868 1352 4924
rect 1352 4868 1356 4924
rect 1292 4864 1356 4868
rect 1372 4924 1436 4928
rect 1372 4868 1376 4924
rect 1376 4868 1432 4924
rect 1432 4868 1436 4924
rect 1372 4864 1436 4868
rect 1452 4924 1516 4928
rect 1452 4868 1456 4924
rect 1456 4868 1512 4924
rect 1512 4868 1516 4924
rect 1452 4864 1516 4868
rect 2484 4924 2548 4928
rect 2484 4868 2488 4924
rect 2488 4868 2544 4924
rect 2544 4868 2548 4924
rect 2484 4864 2548 4868
rect 2564 4924 2628 4928
rect 2564 4868 2568 4924
rect 2568 4868 2624 4924
rect 2624 4868 2628 4924
rect 2564 4864 2628 4868
rect 2644 4924 2708 4928
rect 2644 4868 2648 4924
rect 2648 4868 2704 4924
rect 2704 4868 2708 4924
rect 2644 4864 2708 4868
rect 2724 4924 2788 4928
rect 2724 4868 2728 4924
rect 2728 4868 2784 4924
rect 2784 4868 2788 4924
rect 2724 4864 2788 4868
rect 576 4380 640 4384
rect 576 4324 580 4380
rect 580 4324 636 4380
rect 636 4324 640 4380
rect 576 4320 640 4324
rect 656 4380 720 4384
rect 656 4324 660 4380
rect 660 4324 716 4380
rect 716 4324 720 4380
rect 656 4320 720 4324
rect 736 4380 800 4384
rect 736 4324 740 4380
rect 740 4324 796 4380
rect 796 4324 800 4380
rect 736 4320 800 4324
rect 816 4380 880 4384
rect 816 4324 820 4380
rect 820 4324 876 4380
rect 876 4324 880 4380
rect 816 4320 880 4324
rect 1848 4380 1912 4384
rect 1848 4324 1852 4380
rect 1852 4324 1908 4380
rect 1908 4324 1912 4380
rect 1848 4320 1912 4324
rect 1928 4380 1992 4384
rect 1928 4324 1932 4380
rect 1932 4324 1988 4380
rect 1988 4324 1992 4380
rect 1928 4320 1992 4324
rect 2008 4380 2072 4384
rect 2008 4324 2012 4380
rect 2012 4324 2068 4380
rect 2068 4324 2072 4380
rect 2008 4320 2072 4324
rect 2088 4380 2152 4384
rect 2088 4324 2092 4380
rect 2092 4324 2148 4380
rect 2148 4324 2152 4380
rect 2088 4320 2152 4324
rect 3120 4380 3184 4384
rect 3120 4324 3124 4380
rect 3124 4324 3180 4380
rect 3180 4324 3184 4380
rect 3120 4320 3184 4324
rect 3200 4380 3264 4384
rect 3200 4324 3204 4380
rect 3204 4324 3260 4380
rect 3260 4324 3264 4380
rect 3200 4320 3264 4324
rect 3280 4380 3344 4384
rect 3280 4324 3284 4380
rect 3284 4324 3340 4380
rect 3340 4324 3344 4380
rect 3280 4320 3344 4324
rect 3360 4380 3424 4384
rect 3360 4324 3364 4380
rect 3364 4324 3420 4380
rect 3420 4324 3424 4380
rect 3360 4320 3424 4324
rect 1212 3836 1276 3840
rect 1212 3780 1216 3836
rect 1216 3780 1272 3836
rect 1272 3780 1276 3836
rect 1212 3776 1276 3780
rect 1292 3836 1356 3840
rect 1292 3780 1296 3836
rect 1296 3780 1352 3836
rect 1352 3780 1356 3836
rect 1292 3776 1356 3780
rect 1372 3836 1436 3840
rect 1372 3780 1376 3836
rect 1376 3780 1432 3836
rect 1432 3780 1436 3836
rect 1372 3776 1436 3780
rect 1452 3836 1516 3840
rect 1452 3780 1456 3836
rect 1456 3780 1512 3836
rect 1512 3780 1516 3836
rect 1452 3776 1516 3780
rect 2484 3836 2548 3840
rect 2484 3780 2488 3836
rect 2488 3780 2544 3836
rect 2544 3780 2548 3836
rect 2484 3776 2548 3780
rect 2564 3836 2628 3840
rect 2564 3780 2568 3836
rect 2568 3780 2624 3836
rect 2624 3780 2628 3836
rect 2564 3776 2628 3780
rect 2644 3836 2708 3840
rect 2644 3780 2648 3836
rect 2648 3780 2704 3836
rect 2704 3780 2708 3836
rect 2644 3776 2708 3780
rect 2724 3836 2788 3840
rect 2724 3780 2728 3836
rect 2728 3780 2784 3836
rect 2784 3780 2788 3836
rect 2724 3776 2788 3780
rect 576 3292 640 3296
rect 576 3236 580 3292
rect 580 3236 636 3292
rect 636 3236 640 3292
rect 576 3232 640 3236
rect 656 3292 720 3296
rect 656 3236 660 3292
rect 660 3236 716 3292
rect 716 3236 720 3292
rect 656 3232 720 3236
rect 736 3292 800 3296
rect 736 3236 740 3292
rect 740 3236 796 3292
rect 796 3236 800 3292
rect 736 3232 800 3236
rect 816 3292 880 3296
rect 816 3236 820 3292
rect 820 3236 876 3292
rect 876 3236 880 3292
rect 816 3232 880 3236
rect 1848 3292 1912 3296
rect 1848 3236 1852 3292
rect 1852 3236 1908 3292
rect 1908 3236 1912 3292
rect 1848 3232 1912 3236
rect 1928 3292 1992 3296
rect 1928 3236 1932 3292
rect 1932 3236 1988 3292
rect 1988 3236 1992 3292
rect 1928 3232 1992 3236
rect 2008 3292 2072 3296
rect 2008 3236 2012 3292
rect 2012 3236 2068 3292
rect 2068 3236 2072 3292
rect 2008 3232 2072 3236
rect 2088 3292 2152 3296
rect 2088 3236 2092 3292
rect 2092 3236 2148 3292
rect 2148 3236 2152 3292
rect 2088 3232 2152 3236
rect 3120 3292 3184 3296
rect 3120 3236 3124 3292
rect 3124 3236 3180 3292
rect 3180 3236 3184 3292
rect 3120 3232 3184 3236
rect 3200 3292 3264 3296
rect 3200 3236 3204 3292
rect 3204 3236 3260 3292
rect 3260 3236 3264 3292
rect 3200 3232 3264 3236
rect 3280 3292 3344 3296
rect 3280 3236 3284 3292
rect 3284 3236 3340 3292
rect 3340 3236 3344 3292
rect 3280 3232 3344 3236
rect 3360 3292 3424 3296
rect 3360 3236 3364 3292
rect 3364 3236 3420 3292
rect 3420 3236 3424 3292
rect 3360 3232 3424 3236
rect 1212 2748 1276 2752
rect 1212 2692 1216 2748
rect 1216 2692 1272 2748
rect 1272 2692 1276 2748
rect 1212 2688 1276 2692
rect 1292 2748 1356 2752
rect 1292 2692 1296 2748
rect 1296 2692 1352 2748
rect 1352 2692 1356 2748
rect 1292 2688 1356 2692
rect 1372 2748 1436 2752
rect 1372 2692 1376 2748
rect 1376 2692 1432 2748
rect 1432 2692 1436 2748
rect 1372 2688 1436 2692
rect 1452 2748 1516 2752
rect 1452 2692 1456 2748
rect 1456 2692 1512 2748
rect 1512 2692 1516 2748
rect 1452 2688 1516 2692
rect 2484 2748 2548 2752
rect 2484 2692 2488 2748
rect 2488 2692 2544 2748
rect 2544 2692 2548 2748
rect 2484 2688 2548 2692
rect 2564 2748 2628 2752
rect 2564 2692 2568 2748
rect 2568 2692 2624 2748
rect 2624 2692 2628 2748
rect 2564 2688 2628 2692
rect 2644 2748 2708 2752
rect 2644 2692 2648 2748
rect 2648 2692 2704 2748
rect 2704 2692 2708 2748
rect 2644 2688 2708 2692
rect 2724 2748 2788 2752
rect 2724 2692 2728 2748
rect 2728 2692 2784 2748
rect 2784 2692 2788 2748
rect 2724 2688 2788 2692
rect 576 2204 640 2208
rect 576 2148 580 2204
rect 580 2148 636 2204
rect 636 2148 640 2204
rect 576 2144 640 2148
rect 656 2204 720 2208
rect 656 2148 660 2204
rect 660 2148 716 2204
rect 716 2148 720 2204
rect 656 2144 720 2148
rect 736 2204 800 2208
rect 736 2148 740 2204
rect 740 2148 796 2204
rect 796 2148 800 2204
rect 736 2144 800 2148
rect 816 2204 880 2208
rect 816 2148 820 2204
rect 820 2148 876 2204
rect 876 2148 880 2204
rect 816 2144 880 2148
rect 1848 2204 1912 2208
rect 1848 2148 1852 2204
rect 1852 2148 1908 2204
rect 1908 2148 1912 2204
rect 1848 2144 1912 2148
rect 1928 2204 1992 2208
rect 1928 2148 1932 2204
rect 1932 2148 1988 2204
rect 1988 2148 1992 2204
rect 1928 2144 1992 2148
rect 2008 2204 2072 2208
rect 2008 2148 2012 2204
rect 2012 2148 2068 2204
rect 2068 2148 2072 2204
rect 2008 2144 2072 2148
rect 2088 2204 2152 2208
rect 2088 2148 2092 2204
rect 2092 2148 2148 2204
rect 2148 2148 2152 2204
rect 2088 2144 2152 2148
rect 3120 2204 3184 2208
rect 3120 2148 3124 2204
rect 3124 2148 3180 2204
rect 3180 2148 3184 2204
rect 3120 2144 3184 2148
rect 3200 2204 3264 2208
rect 3200 2148 3204 2204
rect 3204 2148 3260 2204
rect 3260 2148 3264 2204
rect 3200 2144 3264 2148
rect 3280 2204 3344 2208
rect 3280 2148 3284 2204
rect 3284 2148 3340 2204
rect 3340 2148 3344 2204
rect 3280 2144 3344 2148
rect 3360 2204 3424 2208
rect 3360 2148 3364 2204
rect 3364 2148 3420 2204
rect 3420 2148 3424 2204
rect 3360 2144 3424 2148
rect 1212 1660 1276 1664
rect 1212 1604 1216 1660
rect 1216 1604 1272 1660
rect 1272 1604 1276 1660
rect 1212 1600 1276 1604
rect 1292 1660 1356 1664
rect 1292 1604 1296 1660
rect 1296 1604 1352 1660
rect 1352 1604 1356 1660
rect 1292 1600 1356 1604
rect 1372 1660 1436 1664
rect 1372 1604 1376 1660
rect 1376 1604 1432 1660
rect 1432 1604 1436 1660
rect 1372 1600 1436 1604
rect 1452 1660 1516 1664
rect 1452 1604 1456 1660
rect 1456 1604 1512 1660
rect 1512 1604 1516 1660
rect 1452 1600 1516 1604
rect 2484 1660 2548 1664
rect 2484 1604 2488 1660
rect 2488 1604 2544 1660
rect 2544 1604 2548 1660
rect 2484 1600 2548 1604
rect 2564 1660 2628 1664
rect 2564 1604 2568 1660
rect 2568 1604 2624 1660
rect 2624 1604 2628 1660
rect 2564 1600 2628 1604
rect 2644 1660 2708 1664
rect 2644 1604 2648 1660
rect 2648 1604 2704 1660
rect 2704 1604 2708 1660
rect 2644 1600 2708 1604
rect 2724 1660 2788 1664
rect 2724 1604 2728 1660
rect 2728 1604 2784 1660
rect 2784 1604 2788 1660
rect 2724 1600 2788 1604
rect 576 1116 640 1120
rect 576 1060 580 1116
rect 580 1060 636 1116
rect 636 1060 640 1116
rect 576 1056 640 1060
rect 656 1116 720 1120
rect 656 1060 660 1116
rect 660 1060 716 1116
rect 716 1060 720 1116
rect 656 1056 720 1060
rect 736 1116 800 1120
rect 736 1060 740 1116
rect 740 1060 796 1116
rect 796 1060 800 1116
rect 736 1056 800 1060
rect 816 1116 880 1120
rect 816 1060 820 1116
rect 820 1060 876 1116
rect 876 1060 880 1116
rect 816 1056 880 1060
rect 1848 1116 1912 1120
rect 1848 1060 1852 1116
rect 1852 1060 1908 1116
rect 1908 1060 1912 1116
rect 1848 1056 1912 1060
rect 1928 1116 1992 1120
rect 1928 1060 1932 1116
rect 1932 1060 1988 1116
rect 1988 1060 1992 1116
rect 1928 1056 1992 1060
rect 2008 1116 2072 1120
rect 2008 1060 2012 1116
rect 2012 1060 2068 1116
rect 2068 1060 2072 1116
rect 2008 1056 2072 1060
rect 2088 1116 2152 1120
rect 2088 1060 2092 1116
rect 2092 1060 2148 1116
rect 2148 1060 2152 1116
rect 2088 1056 2152 1060
rect 3120 1116 3184 1120
rect 3120 1060 3124 1116
rect 3124 1060 3180 1116
rect 3180 1060 3184 1116
rect 3120 1056 3184 1060
rect 3200 1116 3264 1120
rect 3200 1060 3204 1116
rect 3204 1060 3260 1116
rect 3260 1060 3264 1116
rect 3200 1056 3264 1060
rect 3280 1116 3344 1120
rect 3280 1060 3284 1116
rect 3284 1060 3340 1116
rect 3340 1060 3344 1116
rect 3280 1056 3344 1060
rect 3360 1116 3424 1120
rect 3360 1060 3364 1116
rect 3364 1060 3420 1116
rect 3420 1060 3424 1116
rect 3360 1056 3424 1060
rect 1212 572 1276 576
rect 1212 516 1216 572
rect 1216 516 1272 572
rect 1272 516 1276 572
rect 1212 512 1276 516
rect 1292 572 1356 576
rect 1292 516 1296 572
rect 1296 516 1352 572
rect 1352 516 1356 572
rect 1292 512 1356 516
rect 1372 572 1436 576
rect 1372 516 1376 572
rect 1376 516 1432 572
rect 1432 516 1436 572
rect 1372 512 1436 516
rect 1452 572 1516 576
rect 1452 516 1456 572
rect 1456 516 1512 572
rect 1512 516 1516 572
rect 1452 512 1516 516
rect 2484 572 2548 576
rect 2484 516 2488 572
rect 2488 516 2544 572
rect 2544 516 2548 572
rect 2484 512 2548 516
rect 2564 572 2628 576
rect 2564 516 2568 572
rect 2568 516 2624 572
rect 2624 516 2628 572
rect 2564 512 2628 516
rect 2644 572 2708 576
rect 2644 516 2648 572
rect 2648 516 2704 572
rect 2704 516 2708 572
rect 2644 512 2708 516
rect 2724 572 2788 576
rect 2724 516 2728 572
rect 2728 516 2784 572
rect 2784 516 2788 572
rect 2724 512 2788 516
<< metal4 >>
rect 568 6560 888 7120
rect 568 6496 576 6560
rect 640 6496 656 6560
rect 720 6496 736 6560
rect 800 6496 816 6560
rect 880 6496 888 6560
rect 568 6374 888 6496
rect 568 6138 610 6374
rect 846 6138 888 6374
rect 568 5472 888 6138
rect 568 5408 576 5472
rect 640 5408 656 5472
rect 720 5408 736 5472
rect 800 5408 816 5472
rect 880 5408 888 5472
rect 568 4384 888 5408
rect 568 4320 576 4384
rect 640 4320 656 4384
rect 720 4320 736 4384
rect 800 4320 816 4384
rect 880 4320 888 4384
rect 568 4070 888 4320
rect 568 3834 610 4070
rect 846 3834 888 4070
rect 568 3296 888 3834
rect 568 3232 576 3296
rect 640 3232 656 3296
rect 720 3232 736 3296
rect 800 3232 816 3296
rect 880 3232 888 3296
rect 568 2208 888 3232
rect 568 2144 576 2208
rect 640 2144 656 2208
rect 720 2144 736 2208
rect 800 2144 816 2208
rect 880 2144 888 2208
rect 568 1766 888 2144
rect 568 1530 610 1766
rect 846 1530 888 1766
rect 568 1120 888 1530
rect 568 1056 576 1120
rect 640 1056 656 1120
rect 720 1056 736 1120
rect 800 1056 816 1120
rect 880 1056 888 1120
rect 568 496 888 1056
rect 1204 7104 1524 7120
rect 1204 7040 1212 7104
rect 1276 7040 1292 7104
rect 1356 7040 1372 7104
rect 1436 7040 1452 7104
rect 1516 7040 1524 7104
rect 1204 6016 1524 7040
rect 1204 5952 1212 6016
rect 1276 5952 1292 6016
rect 1356 5952 1372 6016
rect 1436 5952 1452 6016
rect 1516 5952 1524 6016
rect 1204 5222 1524 5952
rect 1204 4986 1246 5222
rect 1482 4986 1524 5222
rect 1204 4928 1524 4986
rect 1204 4864 1212 4928
rect 1276 4864 1292 4928
rect 1356 4864 1372 4928
rect 1436 4864 1452 4928
rect 1516 4864 1524 4928
rect 1204 3840 1524 4864
rect 1204 3776 1212 3840
rect 1276 3776 1292 3840
rect 1356 3776 1372 3840
rect 1436 3776 1452 3840
rect 1516 3776 1524 3840
rect 1204 2918 1524 3776
rect 1204 2752 1246 2918
rect 1482 2752 1524 2918
rect 1204 2688 1212 2752
rect 1516 2688 1524 2752
rect 1204 2682 1246 2688
rect 1482 2682 1524 2688
rect 1204 1664 1524 2682
rect 1204 1600 1212 1664
rect 1276 1600 1292 1664
rect 1356 1600 1372 1664
rect 1436 1600 1452 1664
rect 1516 1600 1524 1664
rect 1204 576 1524 1600
rect 1204 512 1212 576
rect 1276 512 1292 576
rect 1356 512 1372 576
rect 1436 512 1452 576
rect 1516 512 1524 576
rect 1204 496 1524 512
rect 1840 6560 2160 7120
rect 1840 6496 1848 6560
rect 1912 6496 1928 6560
rect 1992 6496 2008 6560
rect 2072 6496 2088 6560
rect 2152 6496 2160 6560
rect 1840 6374 2160 6496
rect 1840 6138 1882 6374
rect 2118 6138 2160 6374
rect 1840 5472 2160 6138
rect 1840 5408 1848 5472
rect 1912 5408 1928 5472
rect 1992 5408 2008 5472
rect 2072 5408 2088 5472
rect 2152 5408 2160 5472
rect 1840 4384 2160 5408
rect 1840 4320 1848 4384
rect 1912 4320 1928 4384
rect 1992 4320 2008 4384
rect 2072 4320 2088 4384
rect 2152 4320 2160 4384
rect 1840 4070 2160 4320
rect 1840 3834 1882 4070
rect 2118 3834 2160 4070
rect 1840 3296 2160 3834
rect 1840 3232 1848 3296
rect 1912 3232 1928 3296
rect 1992 3232 2008 3296
rect 2072 3232 2088 3296
rect 2152 3232 2160 3296
rect 1840 2208 2160 3232
rect 1840 2144 1848 2208
rect 1912 2144 1928 2208
rect 1992 2144 2008 2208
rect 2072 2144 2088 2208
rect 2152 2144 2160 2208
rect 1840 1766 2160 2144
rect 1840 1530 1882 1766
rect 2118 1530 2160 1766
rect 1840 1120 2160 1530
rect 1840 1056 1848 1120
rect 1912 1056 1928 1120
rect 1992 1056 2008 1120
rect 2072 1056 2088 1120
rect 2152 1056 2160 1120
rect 1840 496 2160 1056
rect 2476 7104 2796 7120
rect 2476 7040 2484 7104
rect 2548 7040 2564 7104
rect 2628 7040 2644 7104
rect 2708 7040 2724 7104
rect 2788 7040 2796 7104
rect 2476 6016 2796 7040
rect 2476 5952 2484 6016
rect 2548 5952 2564 6016
rect 2628 5952 2644 6016
rect 2708 5952 2724 6016
rect 2788 5952 2796 6016
rect 2476 5222 2796 5952
rect 2476 4986 2518 5222
rect 2754 4986 2796 5222
rect 2476 4928 2796 4986
rect 2476 4864 2484 4928
rect 2548 4864 2564 4928
rect 2628 4864 2644 4928
rect 2708 4864 2724 4928
rect 2788 4864 2796 4928
rect 2476 3840 2796 4864
rect 2476 3776 2484 3840
rect 2548 3776 2564 3840
rect 2628 3776 2644 3840
rect 2708 3776 2724 3840
rect 2788 3776 2796 3840
rect 2476 2918 2796 3776
rect 2476 2752 2518 2918
rect 2754 2752 2796 2918
rect 2476 2688 2484 2752
rect 2788 2688 2796 2752
rect 2476 2682 2518 2688
rect 2754 2682 2796 2688
rect 2476 1664 2796 2682
rect 2476 1600 2484 1664
rect 2548 1600 2564 1664
rect 2628 1600 2644 1664
rect 2708 1600 2724 1664
rect 2788 1600 2796 1664
rect 2476 576 2796 1600
rect 2476 512 2484 576
rect 2548 512 2564 576
rect 2628 512 2644 576
rect 2708 512 2724 576
rect 2788 512 2796 576
rect 2476 496 2796 512
rect 3112 6560 3432 7120
rect 3112 6496 3120 6560
rect 3184 6496 3200 6560
rect 3264 6496 3280 6560
rect 3344 6496 3360 6560
rect 3424 6496 3432 6560
rect 3112 6374 3432 6496
rect 3112 6138 3154 6374
rect 3390 6138 3432 6374
rect 3112 5472 3432 6138
rect 3112 5408 3120 5472
rect 3184 5408 3200 5472
rect 3264 5408 3280 5472
rect 3344 5408 3360 5472
rect 3424 5408 3432 5472
rect 3112 4384 3432 5408
rect 3112 4320 3120 4384
rect 3184 4320 3200 4384
rect 3264 4320 3280 4384
rect 3344 4320 3360 4384
rect 3424 4320 3432 4384
rect 3112 4070 3432 4320
rect 3112 3834 3154 4070
rect 3390 3834 3432 4070
rect 3112 3296 3432 3834
rect 3112 3232 3120 3296
rect 3184 3232 3200 3296
rect 3264 3232 3280 3296
rect 3344 3232 3360 3296
rect 3424 3232 3432 3296
rect 3112 2208 3432 3232
rect 3112 2144 3120 2208
rect 3184 2144 3200 2208
rect 3264 2144 3280 2208
rect 3344 2144 3360 2208
rect 3424 2144 3432 2208
rect 3112 1766 3432 2144
rect 3112 1530 3154 1766
rect 3390 1530 3432 1766
rect 3112 1120 3432 1530
rect 3112 1056 3120 1120
rect 3184 1056 3200 1120
rect 3264 1056 3280 1120
rect 3344 1056 3360 1120
rect 3424 1056 3432 1120
rect 3112 496 3432 1056
<< via4 >>
rect 610 6138 846 6374
rect 610 3834 846 4070
rect 610 1530 846 1766
rect 1246 4986 1482 5222
rect 1246 2752 1482 2918
rect 1246 2688 1276 2752
rect 1276 2688 1292 2752
rect 1292 2688 1356 2752
rect 1356 2688 1372 2752
rect 1372 2688 1436 2752
rect 1436 2688 1452 2752
rect 1452 2688 1482 2752
rect 1246 2682 1482 2688
rect 1882 6138 2118 6374
rect 1882 3834 2118 4070
rect 1882 1530 2118 1766
rect 2518 4986 2754 5222
rect 2518 2752 2754 2918
rect 2518 2688 2548 2752
rect 2548 2688 2564 2752
rect 2564 2688 2628 2752
rect 2628 2688 2644 2752
rect 2644 2688 2708 2752
rect 2708 2688 2724 2752
rect 2724 2688 2754 2752
rect 2518 2682 2754 2688
rect 3154 6138 3390 6374
rect 3154 3834 3390 4070
rect 3154 1530 3390 1766
<< metal5 >>
rect 92 6374 3864 6416
rect 92 6138 610 6374
rect 846 6138 1882 6374
rect 2118 6138 3154 6374
rect 3390 6138 3864 6374
rect 92 6096 3864 6138
rect 92 5222 3864 5264
rect 92 4986 1246 5222
rect 1482 4986 2518 5222
rect 2754 4986 3864 5222
rect 92 4944 3864 4986
rect 92 4070 3864 4112
rect 92 3834 610 4070
rect 846 3834 1882 4070
rect 2118 3834 3154 4070
rect 3390 3834 3864 4070
rect 92 3792 3864 3834
rect 92 2918 3864 2960
rect 92 2682 1246 2918
rect 1482 2682 2518 2918
rect 2754 2682 3864 2918
rect 92 2640 3864 2682
rect 92 1766 3864 1808
rect 92 1530 610 1766
rect 846 1530 1882 1766
rect 2118 1530 3154 1766
rect 3390 1530 3864 1766
rect 92 1488 3864 1530
use sky130_fd_sc_hd__and3b_1  _07_
timestamp 1694031861
transform -1 0 1932 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _08_
timestamp 1694031861
transform -1 0 1012 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _09_
timestamp 1694031861
transform 1 0 2300 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  _10_
timestamp 1694031861
transform 1 0 1932 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  _11_
timestamp 1694031861
transform -1 0 1472 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__nor3b_2  _12_
timestamp 1694031861
transform -1 0 1840 0 -1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__nor3b_2  _13_
timestamp 1694031861
transform -1 0 2852 0 -1 3808
box -38 -48 958 592
use sky130_fd_sc_hd__nor3_2  _14_
timestamp 1694031861
transform -1 0 2944 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__nor3b_2  _15_
timestamp 1694031861
transform 1 0 1104 0 1 1632
box -38 -48 958 592
use sky130_fd_sc_hd__and3b_1  _16_
timestamp 1694031861
transform -1 0 2300 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _17_
timestamp 1694031861
transform -1 0 920 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _18_
timestamp 1694031861
transform 1 0 1380 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1694031861
transform -1 0 3036 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _20_
timestamp 1694031861
transform 1 0 368 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1694031861
transform 1 0 1104 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7
timestamp 1694031861
transform 1 0 736 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1694031861
transform 1 0 2300 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29
timestamp 1694031861
transform 1 0 2760 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34
timestamp 1694031861
transform 1 0 3220 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1694031861
transform 1 0 368 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_10
timestamp 1694031861
transform 1 0 1012 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_21
timestamp 1694031861
transform 1 0 2024 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_34
timestamp 1694031861
transform 1 0 3220 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1694031861
transform 1 0 368 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_21
timestamp 1694031861
transform 1 0 2024 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1694031861
transform 1 0 2576 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_32
timestamp 1694031861
transform 1 0 3036 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1694031861
transform 1 0 368 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_9
timestamp 1694031861
transform 1 0 920 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_20
timestamp 1694031861
transform 1 0 1932 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_33
timestamp 1694031861
transform 1 0 3128 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_37
timestamp 1694031861
transform 1 0 3496 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1694031861
transform 1 0 368 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_13
timestamp 1694031861
transform 1 0 1288 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1694031861
transform 1 0 2300 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_29
timestamp 1694031861
transform 1 0 2760 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_37
timestamp 1694031861
transform 1 0 3496 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_12
timestamp 1694031861
transform 1 0 1196 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_30
timestamp 1694031861
transform 1 0 2852 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1694031861
transform 1 0 368 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1694031861
transform 1 0 1472 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1694031861
transform 1 0 2576 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_29
timestamp 1694031861
transform 1 0 2760 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_34
timestamp 1694031861
transform 1 0 3220 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1694031861
transform 1 0 368 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_19
timestamp 1694031861
transform 1 0 1840 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_31
timestamp 1694031861
transform 1 0 2944 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_37
timestamp 1694031861
transform 1 0 3496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_8
timestamp 1694031861
transform 1 0 828 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_16
timestamp 1694031861
transform 1 0 1564 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1694031861
transform 1 0 2300 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_29
timestamp 1694031861
transform 1 0 2760 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_37
timestamp 1694031861
transform 1 0 3496 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1694031861
transform 1 0 368 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_15
timestamp 1694031861
transform 1 0 1472 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_19
timestamp 1694031861
transform 1 0 1840 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_29
timestamp 1694031861
transform 1 0 2760 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_37
timestamp 1694031861
transform 1 0 3496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1694031861
transform 1 0 368 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_15
timestamp 1694031861
transform 1 0 1472 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1694031861
transform 1 0 2300 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_29
timestamp 1694031861
transform 1 0 2760 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_37
timestamp 1694031861
transform 1 0 3496 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_12
timestamp 1694031861
transform 1 0 1196 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_24
timestamp 1694031861
transform 1 0 2300 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_29
timestamp 1694031861
transform 1 0 2760 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_37
timestamp 1694031861
transform 1 0 3496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_6  input1
timestamp 1694031861
transform 1 0 368 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  input2
timestamp 1694031861
transform 1 0 368 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1694031861
transform 1 0 368 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output4
timestamp 1694031861
transform -1 0 2300 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output5
timestamp 1694031861
transform -1 0 2300 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  output6
timestamp 1694031861
transform 1 0 1748 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1694031861
transform 1 0 2852 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output8
timestamp 1694031861
transform -1 0 1288 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  output9
timestamp 1694031861
transform 1 0 2392 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1694031861
transform 1 0 2852 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  output11
timestamp 1694031861
transform 1 0 1472 0 1 544
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1694031861
transform 1 0 92 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1694031861
transform -1 0 3864 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1694031861
transform 1 0 92 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1694031861
transform -1 0 3864 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1694031861
transform 1 0 92 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1694031861
transform -1 0 3864 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1694031861
transform 1 0 92 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1694031861
transform -1 0 3864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1694031861
transform 1 0 92 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1694031861
transform -1 0 3864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1694031861
transform 1 0 92 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1694031861
transform -1 0 3864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1694031861
transform 1 0 92 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1694031861
transform -1 0 3864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1694031861
transform 1 0 92 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1694031861
transform -1 0 3864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1694031861
transform 1 0 92 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1694031861
transform -1 0 3864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1694031861
transform 1 0 92 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1694031861
transform -1 0 3864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1694031861
transform 1 0 92 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1694031861
transform -1 0 3864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1694031861
transform 1 0 92 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1694031861
transform -1 0 3864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1694031861
transform 1 0 2668 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1694031861
transform 1 0 2668 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1694031861
transform 1 0 2668 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1694031861
transform 1 0 2668 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1694031861
transform 1 0 2668 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1694031861
transform 1 0 2668 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1694031861
transform 1 0 2668 0 -1 7072
box -38 -48 130 592
<< labels >>
rlabel metal3 s 0 6566 200 6626 4 in[0]
port 1 nsew
rlabel metal3 s 0 3846 200 3906 4 in[1]
port 2 nsew
rlabel metal3 s 0 1262 200 1322 4 in[2]
port 3 nsew
rlabel metal3 s 3800 7182 4000 7242 4 out[0]
port 4 nsew
rlabel metal3 s 3800 6430 4000 6490 4 out[1]
port 5 nsew
rlabel metal3 s 3800 5342 4000 5402 4 out[2]
port 6 nsew
rlabel metal3 s 3800 4390 4000 4450 4 out[3]
port 7 nsew
rlabel metal3 s 3800 3438 4000 3498 4 out[4]
port 8 nsew
rlabel metal3 s 3800 2350 4000 2410 4 out[5]
port 9 nsew
rlabel metal3 s 3800 1398 4000 1458 4 out[6]
port 10 nsew
rlabel metal3 s 3800 446 4000 506 4 out[7]
port 11 nsew
rlabel metal4 s 1204 496 1524 7120 4 VGND
port 12 nsew
rlabel metal4 s 2476 496 2796 7120 4 VGND
port 12 nsew
rlabel metal5 s 92 2640 3864 2960 4 VGND
port 12 nsew
rlabel metal5 s 92 4944 3864 5264 4 VGND
port 12 nsew
rlabel metal4 s 568 496 888 7120 4 VPWR
port 13 nsew
rlabel metal4 s 1840 496 2160 7120 4 VPWR
port 13 nsew
rlabel metal4 s 3112 496 3432 7120 4 VPWR
port 13 nsew
rlabel metal5 s 92 1488 3864 1808 4 VPWR
port 13 nsew
rlabel metal5 s 92 3792 3864 4112 4 VPWR
port 13 nsew
rlabel metal5 s 92 6096 3864 6416 4 VPWR
port 13 nsew
<< properties >>
string FIXED_BBOX 0 0 4000 8000
<< end >>
