magic
tech sky130A
timestamp 1699926577
<< metal1 >>
rect -5 586 97 601
rect -5 16 17 586
rect 75 16 97 586
rect -5 1 97 16
<< via1 >>
rect 17 16 75 586
<< metal2 >>
rect -7 586 98 600
rect -7 575 17 586
rect 75 575 98 586
rect -7 27 12 575
rect 80 27 98 575
rect -7 16 17 27
rect 75 16 98 27
rect -7 -2 98 16
<< via2 >>
rect 12 27 17 575
rect 17 27 75 575
rect 75 27 80 575
<< metal3 >>
rect -7 577 98 600
rect -7 575 30 577
rect 62 575 98 577
rect -7 27 12 575
rect 80 27 98 575
rect -7 25 30 27
rect 62 25 98 27
rect -7 -2 98 25
<< via3 >>
rect 30 575 62 577
rect 30 545 62 575
rect 30 505 62 537
rect 30 465 62 497
rect 30 425 62 457
rect 30 385 62 417
rect 30 345 62 377
rect 30 305 62 337
rect 30 265 62 297
rect 30 225 62 257
rect 30 185 62 217
rect 30 145 62 177
rect 30 105 62 137
rect 30 65 62 97
rect 30 27 62 57
rect 30 25 62 27
<< metal4 >>
rect -7 577 98 600
rect -7 545 30 577
rect 62 545 98 577
rect -7 537 98 545
rect -7 505 30 537
rect 62 505 98 537
rect -7 497 98 505
rect -7 465 30 497
rect 62 465 98 497
rect -7 457 98 465
rect -7 425 30 457
rect 62 425 98 457
rect -7 417 98 425
rect -7 385 30 417
rect 62 385 98 417
rect -7 377 98 385
rect -7 345 30 377
rect 62 345 98 377
rect -7 337 98 345
rect -7 305 30 337
rect 62 305 98 337
rect -7 297 98 305
rect -7 265 30 297
rect 62 265 98 297
rect -7 257 98 265
rect -7 225 30 257
rect 62 225 98 257
rect -7 217 98 225
rect -7 185 30 217
rect 62 185 98 217
rect -7 177 98 185
rect -7 145 30 177
rect 62 145 98 177
rect -7 137 98 145
rect -7 105 30 137
rect 62 105 98 137
rect -7 97 98 105
rect -7 65 30 97
rect 62 65 98 97
rect -7 57 98 65
rect -7 25 30 57
rect 62 25 98 57
rect -7 -2 98 25
<< end >>
