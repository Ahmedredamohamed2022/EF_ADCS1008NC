magic
tech sky130A
magscale 1 2
timestamp 1699926577
<< metal3 >>
rect -1186 2312 1186 2340
rect -1186 2248 1102 2312
rect 1166 2248 1186 2312
rect -1186 2232 1186 2248
rect -1186 2168 1102 2232
rect 1166 2168 1186 2232
rect -1186 2152 1186 2168
rect -1186 2088 1102 2152
rect 1166 2088 1186 2152
rect -1186 2072 1186 2088
rect -1186 2008 1102 2072
rect 1166 2008 1186 2072
rect -1186 1992 1186 2008
rect -1186 1928 1102 1992
rect 1166 1928 1186 1992
rect -1186 1912 1186 1928
rect -1186 1848 1102 1912
rect 1166 1848 1186 1912
rect -1186 1832 1186 1848
rect -1186 1768 1102 1832
rect 1166 1768 1186 1832
rect -1186 1752 1186 1768
rect -1186 1688 1102 1752
rect 1166 1688 1186 1752
rect -1186 1672 1186 1688
rect -1186 1608 1102 1672
rect 1166 1608 1186 1672
rect -1186 1592 1186 1608
rect -1186 1528 1102 1592
rect 1166 1528 1186 1592
rect -1186 1512 1186 1528
rect -1186 1448 1102 1512
rect 1166 1448 1186 1512
rect -1186 1432 1186 1448
rect -1186 1368 1102 1432
rect 1166 1368 1186 1432
rect -1186 1352 1186 1368
rect -1186 1288 1102 1352
rect 1166 1288 1186 1352
rect -1186 1272 1186 1288
rect -1186 1208 1102 1272
rect 1166 1208 1186 1272
rect -1186 1192 1186 1208
rect -1186 1128 1102 1192
rect 1166 1128 1186 1192
rect -1186 1112 1186 1128
rect -1186 1048 1102 1112
rect 1166 1048 1186 1112
rect -1186 1032 1186 1048
rect -1186 968 1102 1032
rect 1166 968 1186 1032
rect -1186 952 1186 968
rect -1186 888 1102 952
rect 1166 888 1186 952
rect -1186 872 1186 888
rect -1186 808 1102 872
rect 1166 808 1186 872
rect -1186 792 1186 808
rect -1186 728 1102 792
rect 1166 728 1186 792
rect -1186 712 1186 728
rect -1186 648 1102 712
rect 1166 648 1186 712
rect -1186 632 1186 648
rect -1186 568 1102 632
rect 1166 568 1186 632
rect -1186 552 1186 568
rect -1186 488 1102 552
rect 1166 488 1186 552
rect -1186 472 1186 488
rect -1186 408 1102 472
rect 1166 408 1186 472
rect -1186 392 1186 408
rect -1186 328 1102 392
rect 1166 328 1186 392
rect -1186 312 1186 328
rect -1186 248 1102 312
rect 1166 248 1186 312
rect -1186 232 1186 248
rect -1186 168 1102 232
rect 1166 168 1186 232
rect -1186 152 1186 168
rect -1186 88 1102 152
rect 1166 88 1186 152
rect -1186 72 1186 88
rect -1186 8 1102 72
rect 1166 8 1186 72
rect -1186 -8 1186 8
rect -1186 -72 1102 -8
rect 1166 -72 1186 -8
rect -1186 -88 1186 -72
rect -1186 -152 1102 -88
rect 1166 -152 1186 -88
rect -1186 -168 1186 -152
rect -1186 -232 1102 -168
rect 1166 -232 1186 -168
rect -1186 -248 1186 -232
rect -1186 -312 1102 -248
rect 1166 -312 1186 -248
rect -1186 -328 1186 -312
rect -1186 -392 1102 -328
rect 1166 -392 1186 -328
rect -1186 -408 1186 -392
rect -1186 -472 1102 -408
rect 1166 -472 1186 -408
rect -1186 -488 1186 -472
rect -1186 -552 1102 -488
rect 1166 -552 1186 -488
rect -1186 -568 1186 -552
rect -1186 -632 1102 -568
rect 1166 -632 1186 -568
rect -1186 -648 1186 -632
rect -1186 -712 1102 -648
rect 1166 -712 1186 -648
rect -1186 -728 1186 -712
rect -1186 -792 1102 -728
rect 1166 -792 1186 -728
rect -1186 -808 1186 -792
rect -1186 -872 1102 -808
rect 1166 -872 1186 -808
rect -1186 -888 1186 -872
rect -1186 -952 1102 -888
rect 1166 -952 1186 -888
rect -1186 -968 1186 -952
rect -1186 -1032 1102 -968
rect 1166 -1032 1186 -968
rect -1186 -1048 1186 -1032
rect -1186 -1112 1102 -1048
rect 1166 -1112 1186 -1048
rect -1186 -1128 1186 -1112
rect -1186 -1192 1102 -1128
rect 1166 -1192 1186 -1128
rect -1186 -1208 1186 -1192
rect -1186 -1272 1102 -1208
rect 1166 -1272 1186 -1208
rect -1186 -1288 1186 -1272
rect -1186 -1352 1102 -1288
rect 1166 -1352 1186 -1288
rect -1186 -1368 1186 -1352
rect -1186 -1432 1102 -1368
rect 1166 -1432 1186 -1368
rect -1186 -1448 1186 -1432
rect -1186 -1512 1102 -1448
rect 1166 -1512 1186 -1448
rect -1186 -1528 1186 -1512
rect -1186 -1592 1102 -1528
rect 1166 -1592 1186 -1528
rect -1186 -1608 1186 -1592
rect -1186 -1672 1102 -1608
rect 1166 -1672 1186 -1608
rect -1186 -1688 1186 -1672
rect -1186 -1752 1102 -1688
rect 1166 -1752 1186 -1688
rect -1186 -1768 1186 -1752
rect -1186 -1832 1102 -1768
rect 1166 -1832 1186 -1768
rect -1186 -1848 1186 -1832
rect -1186 -1912 1102 -1848
rect 1166 -1912 1186 -1848
rect -1186 -1928 1186 -1912
rect -1186 -1992 1102 -1928
rect 1166 -1992 1186 -1928
rect -1186 -2008 1186 -1992
rect -1186 -2072 1102 -2008
rect 1166 -2072 1186 -2008
rect -1186 -2088 1186 -2072
rect -1186 -2152 1102 -2088
rect 1166 -2152 1186 -2088
rect -1186 -2168 1186 -2152
rect -1186 -2232 1102 -2168
rect 1166 -2232 1186 -2168
rect -1186 -2248 1186 -2232
rect -1186 -2312 1102 -2248
rect 1166 -2312 1186 -2248
rect -1186 -2340 1186 -2312
<< via3 >>
rect 1102 2248 1166 2312
rect 1102 2168 1166 2232
rect 1102 2088 1166 2152
rect 1102 2008 1166 2072
rect 1102 1928 1166 1992
rect 1102 1848 1166 1912
rect 1102 1768 1166 1832
rect 1102 1688 1166 1752
rect 1102 1608 1166 1672
rect 1102 1528 1166 1592
rect 1102 1448 1166 1512
rect 1102 1368 1166 1432
rect 1102 1288 1166 1352
rect 1102 1208 1166 1272
rect 1102 1128 1166 1192
rect 1102 1048 1166 1112
rect 1102 968 1166 1032
rect 1102 888 1166 952
rect 1102 808 1166 872
rect 1102 728 1166 792
rect 1102 648 1166 712
rect 1102 568 1166 632
rect 1102 488 1166 552
rect 1102 408 1166 472
rect 1102 328 1166 392
rect 1102 248 1166 312
rect 1102 168 1166 232
rect 1102 88 1166 152
rect 1102 8 1166 72
rect 1102 -72 1166 -8
rect 1102 -152 1166 -88
rect 1102 -232 1166 -168
rect 1102 -312 1166 -248
rect 1102 -392 1166 -328
rect 1102 -472 1166 -408
rect 1102 -552 1166 -488
rect 1102 -632 1166 -568
rect 1102 -712 1166 -648
rect 1102 -792 1166 -728
rect 1102 -872 1166 -808
rect 1102 -952 1166 -888
rect 1102 -1032 1166 -968
rect 1102 -1112 1166 -1048
rect 1102 -1192 1166 -1128
rect 1102 -1272 1166 -1208
rect 1102 -1352 1166 -1288
rect 1102 -1432 1166 -1368
rect 1102 -1512 1166 -1448
rect 1102 -1592 1166 -1528
rect 1102 -1672 1166 -1608
rect 1102 -1752 1166 -1688
rect 1102 -1832 1166 -1768
rect 1102 -1912 1166 -1848
rect 1102 -1992 1166 -1928
rect 1102 -2072 1166 -2008
rect 1102 -2152 1166 -2088
rect 1102 -2232 1166 -2168
rect 1102 -2312 1166 -2248
<< mimcap >>
rect -1146 2232 854 2300
rect -1146 -2232 -1098 2232
rect 806 -2232 854 2232
rect -1146 -2300 854 -2232
<< mimcapcontact >>
rect -1098 -2232 806 2232
<< metal4 >>
rect 1086 2312 1182 2328
rect -1107 2232 815 2261
rect -1107 -2232 -1098 2232
rect 806 -2232 815 2232
rect -1107 -2261 815 -2232
rect 1086 2248 1102 2312
rect 1166 2248 1182 2312
rect 1086 2232 1182 2248
rect 1086 2168 1102 2232
rect 1166 2168 1182 2232
rect 1086 2152 1182 2168
rect 1086 2088 1102 2152
rect 1166 2088 1182 2152
rect 1086 2072 1182 2088
rect 1086 2008 1102 2072
rect 1166 2008 1182 2072
rect 1086 1992 1182 2008
rect 1086 1928 1102 1992
rect 1166 1928 1182 1992
rect 1086 1912 1182 1928
rect 1086 1848 1102 1912
rect 1166 1848 1182 1912
rect 1086 1832 1182 1848
rect 1086 1768 1102 1832
rect 1166 1768 1182 1832
rect 1086 1752 1182 1768
rect 1086 1688 1102 1752
rect 1166 1688 1182 1752
rect 1086 1672 1182 1688
rect 1086 1608 1102 1672
rect 1166 1608 1182 1672
rect 1086 1592 1182 1608
rect 1086 1528 1102 1592
rect 1166 1528 1182 1592
rect 1086 1512 1182 1528
rect 1086 1448 1102 1512
rect 1166 1448 1182 1512
rect 1086 1432 1182 1448
rect 1086 1368 1102 1432
rect 1166 1368 1182 1432
rect 1086 1352 1182 1368
rect 1086 1288 1102 1352
rect 1166 1288 1182 1352
rect 1086 1272 1182 1288
rect 1086 1208 1102 1272
rect 1166 1208 1182 1272
rect 1086 1192 1182 1208
rect 1086 1128 1102 1192
rect 1166 1128 1182 1192
rect 1086 1112 1182 1128
rect 1086 1048 1102 1112
rect 1166 1048 1182 1112
rect 1086 1032 1182 1048
rect 1086 968 1102 1032
rect 1166 968 1182 1032
rect 1086 952 1182 968
rect 1086 888 1102 952
rect 1166 888 1182 952
rect 1086 872 1182 888
rect 1086 808 1102 872
rect 1166 808 1182 872
rect 1086 792 1182 808
rect 1086 728 1102 792
rect 1166 728 1182 792
rect 1086 712 1182 728
rect 1086 648 1102 712
rect 1166 648 1182 712
rect 1086 632 1182 648
rect 1086 568 1102 632
rect 1166 568 1182 632
rect 1086 552 1182 568
rect 1086 488 1102 552
rect 1166 488 1182 552
rect 1086 472 1182 488
rect 1086 408 1102 472
rect 1166 408 1182 472
rect 1086 392 1182 408
rect 1086 328 1102 392
rect 1166 328 1182 392
rect 1086 312 1182 328
rect 1086 248 1102 312
rect 1166 248 1182 312
rect 1086 232 1182 248
rect 1086 168 1102 232
rect 1166 168 1182 232
rect 1086 152 1182 168
rect 1086 88 1102 152
rect 1166 88 1182 152
rect 1086 72 1182 88
rect 1086 8 1102 72
rect 1166 8 1182 72
rect 1086 -8 1182 8
rect 1086 -72 1102 -8
rect 1166 -72 1182 -8
rect 1086 -88 1182 -72
rect 1086 -152 1102 -88
rect 1166 -152 1182 -88
rect 1086 -168 1182 -152
rect 1086 -232 1102 -168
rect 1166 -232 1182 -168
rect 1086 -248 1182 -232
rect 1086 -312 1102 -248
rect 1166 -312 1182 -248
rect 1086 -328 1182 -312
rect 1086 -392 1102 -328
rect 1166 -392 1182 -328
rect 1086 -408 1182 -392
rect 1086 -472 1102 -408
rect 1166 -472 1182 -408
rect 1086 -488 1182 -472
rect 1086 -552 1102 -488
rect 1166 -552 1182 -488
rect 1086 -568 1182 -552
rect 1086 -632 1102 -568
rect 1166 -632 1182 -568
rect 1086 -648 1182 -632
rect 1086 -712 1102 -648
rect 1166 -712 1182 -648
rect 1086 -728 1182 -712
rect 1086 -792 1102 -728
rect 1166 -792 1182 -728
rect 1086 -808 1182 -792
rect 1086 -872 1102 -808
rect 1166 -872 1182 -808
rect 1086 -888 1182 -872
rect 1086 -952 1102 -888
rect 1166 -952 1182 -888
rect 1086 -968 1182 -952
rect 1086 -1032 1102 -968
rect 1166 -1032 1182 -968
rect 1086 -1048 1182 -1032
rect 1086 -1112 1102 -1048
rect 1166 -1112 1182 -1048
rect 1086 -1128 1182 -1112
rect 1086 -1192 1102 -1128
rect 1166 -1192 1182 -1128
rect 1086 -1208 1182 -1192
rect 1086 -1272 1102 -1208
rect 1166 -1272 1182 -1208
rect 1086 -1288 1182 -1272
rect 1086 -1352 1102 -1288
rect 1166 -1352 1182 -1288
rect 1086 -1368 1182 -1352
rect 1086 -1432 1102 -1368
rect 1166 -1432 1182 -1368
rect 1086 -1448 1182 -1432
rect 1086 -1512 1102 -1448
rect 1166 -1512 1182 -1448
rect 1086 -1528 1182 -1512
rect 1086 -1592 1102 -1528
rect 1166 -1592 1182 -1528
rect 1086 -1608 1182 -1592
rect 1086 -1672 1102 -1608
rect 1166 -1672 1182 -1608
rect 1086 -1688 1182 -1672
rect 1086 -1752 1102 -1688
rect 1166 -1752 1182 -1688
rect 1086 -1768 1182 -1752
rect 1086 -1832 1102 -1768
rect 1166 -1832 1182 -1768
rect 1086 -1848 1182 -1832
rect 1086 -1912 1102 -1848
rect 1166 -1912 1182 -1848
rect 1086 -1928 1182 -1912
rect 1086 -1992 1102 -1928
rect 1166 -1992 1182 -1928
rect 1086 -2008 1182 -1992
rect 1086 -2072 1102 -2008
rect 1166 -2072 1182 -2008
rect 1086 -2088 1182 -2072
rect 1086 -2152 1102 -2088
rect 1166 -2152 1182 -2088
rect 1086 -2168 1182 -2152
rect 1086 -2232 1102 -2168
rect 1166 -2232 1182 -2168
rect 1086 -2248 1182 -2232
rect 1086 -2312 1102 -2248
rect 1166 -2312 1182 -2248
rect 1086 -2328 1182 -2312
<< properties >>
string FIXED_BBOX -1186 -2340 894 2340
<< end >>
