magic
tech sky130A
magscale 1 2
timestamp 1699522684
<< metal1 >>
rect 788 90863 1322 90889
rect 788 90831 801 90863
rect 784 90747 801 90831
rect 1301 90831 1322 90863
rect 1301 90747 2290 90831
rect 784 90727 2290 90747
rect 1806 88021 2212 88046
rect 1806 87777 1823 88021
rect 2195 87777 2212 88021
rect 1806 87752 2212 87777
rect 11 87218 1368 87223
rect 11 87196 1374 87218
rect 11 87080 37 87196
rect 601 87080 1374 87196
rect 11 87021 1374 87080
rect 1174 87018 1374 87021
rect 1420 84540 1702 84564
rect 1420 84296 1439 84540
rect 1683 84296 1702 84540
rect 1420 84272 1702 84296
rect 3016 84080 3316 84126
rect 3016 83452 3048 84080
rect 3292 83452 3316 84080
rect 3016 83392 3316 83452
rect 790 83253 1374 83298
rect 790 83137 825 83253
rect 1325 83137 1374 83253
rect 790 83100 1374 83137
rect 812 83098 1374 83100
rect 34580 82977 35070 82985
rect 1168 82953 1374 82962
rect 806 82919 1450 82953
rect 806 82803 844 82919
rect 1408 82803 1450 82919
rect 33304 82939 35070 82977
rect 21068 82885 21262 82889
rect 806 82769 1450 82803
rect 20506 82846 21262 82885
rect 1168 82752 1374 82769
rect 20506 82730 21109 82846
rect 21225 82730 21262 82846
rect 20506 82687 21262 82730
rect 20510 82686 20642 82687
rect 33304 82631 34639 82939
rect 35011 82631 35070 82939
rect 33304 82569 35070 82631
<< via1 >>
rect 801 90747 1301 90863
rect 1823 87777 2195 88021
rect 37 87080 601 87196
rect 1439 84296 1683 84540
rect 3048 83452 3292 84080
rect 825 83137 1325 83253
rect 844 82803 1408 82919
rect 21109 82730 21225 82846
rect 34639 82631 35011 82939
<< metal2 >>
rect 4424 103475 4520 103773
rect 7828 103473 7918 103773
rect 11230 103465 11320 103773
rect 14528 103465 14618 103773
rect 17840 103467 17936 103773
rect 21214 103467 21310 103773
rect 24516 103467 24612 103773
rect 27962 103465 28050 103773
rect 35196 103719 35256 103773
rect 35342 103719 35402 103773
rect 35488 103721 35548 103773
rect 35188 103681 35268 103719
rect 35188 103625 35203 103681
rect 35259 103625 35268 103681
rect 35188 103585 35268 103625
rect 35336 103685 35412 103719
rect 35336 103629 35346 103685
rect 35402 103629 35412 103685
rect 35336 103585 35412 103629
rect 35480 103683 35556 103721
rect 35480 103627 35494 103683
rect 35550 103627 35556 103683
rect 35480 103585 35556 103627
rect 36404 103599 36598 103773
rect 36404 103383 36426 103599
rect 36562 103383 36598 103599
rect 36404 103333 36598 103383
rect 27882 99499 28140 99555
rect 27882 99281 27899 99499
rect 27870 99043 27899 99281
rect 28115 99043 28140 99499
rect 27870 98981 28140 99043
rect 27870 98783 28132 98981
rect 788 90873 1322 90889
rect 788 90863 823 90873
rect 1279 90863 1322 90873
rect 788 90747 801 90863
rect 1301 90747 1322 90863
rect 788 90737 823 90747
rect 1279 90737 1322 90747
rect 788 90727 1322 90737
rect 1786 90653 2122 90663
rect 1786 90597 1805 90653
rect 1861 90597 1885 90653
rect 1941 90597 1965 90653
rect 2021 90597 2045 90653
rect 2101 90597 2122 90653
rect 1410 90474 1720 90494
rect 1410 90418 1455 90474
rect 1511 90418 1535 90474
rect 1591 90418 1615 90474
rect 1671 90418 1720 90474
rect 1410 88066 1720 90418
rect 1408 87736 1720 88066
rect 2 87206 632 87235
rect 2 87196 51 87206
rect 587 87196 632 87206
rect 2 87080 37 87196
rect 601 87080 632 87196
rect 2 87070 51 87080
rect 587 87070 632 87080
rect 2 87033 632 87070
rect 1410 84540 1720 87736
rect 1786 88382 2122 90597
rect 27910 90479 28132 98783
rect 27910 90423 27950 90479
rect 28006 90423 28030 90479
rect 28086 90423 28132 90479
rect 27910 90402 28132 90423
rect 3012 90287 3312 90331
rect 3012 89991 3053 90287
rect 3269 89991 3312 90287
rect 1786 88068 2240 88382
rect 1786 88021 2246 88068
rect 1786 87777 1823 88021
rect 2195 87777 2246 88021
rect 1786 87718 2246 87777
rect 1410 84296 1439 84540
rect 1683 84296 1720 84540
rect 1410 84267 1720 84296
rect 3012 84126 3312 89991
rect 3012 84080 3316 84126
rect 3012 83452 3048 84080
rect 3292 83452 3316 84080
rect 3012 83418 3316 83452
rect 3016 83392 3316 83418
rect 790 83263 1374 83298
rect 790 83253 847 83263
rect 1303 83253 1374 83263
rect 790 83137 825 83253
rect 1325 83137 1374 83253
rect 790 83127 847 83137
rect 1303 83127 1374 83137
rect 790 83100 1374 83127
rect 806 82929 1450 82953
rect 806 82919 858 82929
rect 1394 82919 1450 82929
rect 806 82803 844 82919
rect 1408 82803 1450 82919
rect 34580 82939 35070 82985
rect 34580 82933 34639 82939
rect 35011 82933 35070 82939
rect 806 82793 858 82803
rect 1394 82793 1450 82803
rect 806 82769 1450 82793
rect 21068 82856 21262 82889
rect 21068 82720 21099 82856
rect 21235 82720 21262 82856
rect 21068 82689 21262 82720
rect 34580 82637 34637 82933
rect 35013 82637 35070 82933
rect 34580 82631 34639 82637
rect 35011 82631 35070 82637
rect 34580 82577 35070 82631
rect 33630 80424 33806 80553
rect 33630 80288 33647 80424
rect 33783 80288 33806 80424
rect 33630 80257 33806 80288
rect 19202 77476 19814 77561
rect 19202 77020 19305 77476
rect 19681 77020 19814 77476
rect 19202 76951 19814 77020
rect 19346 76027 19610 76951
rect 23594 76519 24210 76587
rect 23594 76063 23659 76519
rect 24115 76063 24210 76519
rect 32200 76233 32752 76235
rect 19374 75699 19596 76027
rect 23594 75993 24210 76063
rect 32198 76144 32762 76233
rect 23770 75707 23986 75993
rect 32198 75768 32252 76144
rect 32708 75768 32762 76144
rect 32198 75695 32762 75768
rect 32200 75677 32752 75695
rect 32336 75577 32558 75677
<< via2 >>
rect 35203 103625 35259 103681
rect 35346 103629 35402 103685
rect 35494 103627 35550 103683
rect 36426 103383 36562 103599
rect 27899 99043 28115 99499
rect 823 90863 1279 90873
rect 823 90747 1279 90863
rect 823 90737 1279 90747
rect 1805 90597 1861 90653
rect 1885 90597 1941 90653
rect 1965 90597 2021 90653
rect 2045 90597 2101 90653
rect 1455 90418 1511 90474
rect 1535 90418 1591 90474
rect 1615 90418 1671 90474
rect 51 87196 587 87206
rect 51 87080 587 87196
rect 51 87070 587 87080
rect 27950 90423 28006 90479
rect 28030 90423 28086 90479
rect 3053 89991 3269 90287
rect 847 83253 1303 83263
rect 847 83137 1303 83253
rect 847 83127 1303 83137
rect 858 82919 1394 82929
rect 858 82803 1394 82919
rect 858 82793 1394 82803
rect 21099 82846 21235 82856
rect 21099 82730 21109 82846
rect 21109 82730 21225 82846
rect 21225 82730 21235 82846
rect 21099 82720 21235 82730
rect 34637 82637 34639 82933
rect 34639 82637 35011 82933
rect 35011 82637 35013 82933
rect 33647 80288 33783 80424
rect 19305 77020 19681 77476
rect 23659 76063 24115 76519
rect 32252 75768 32708 76144
<< metal3 >>
rect 35341 103719 35402 103743
rect 35488 103721 35548 103743
rect 35188 103681 35268 103719
rect 35188 103625 35203 103681
rect 35259 103625 35268 103681
rect 35188 103585 35268 103625
rect 35336 103685 35412 103719
rect 35336 103629 35346 103685
rect 35402 103629 35412 103685
rect 35336 103585 35412 103629
rect 35480 103683 35556 103721
rect 35480 103627 35494 103683
rect 35550 103627 35556 103683
rect 35480 103585 35556 103627
rect 36406 103599 36598 103653
rect 27882 99503 28140 99555
rect 27882 99039 27895 99503
rect 28119 99039 28140 99503
rect 27882 98981 28140 99039
rect 35196 97643 35256 103585
rect 34802 97583 35256 97643
rect 35341 97505 35402 103585
rect 34910 97445 35402 97505
rect 35107 97444 35402 97445
rect 35107 97443 35363 97444
rect 35488 97371 35548 103585
rect 34812 97311 35548 97371
rect 36406 103383 36426 103599
rect 36562 103383 36598 103599
rect 21304 95045 21512 95085
rect 21304 94981 21335 95045
rect 21399 94981 21415 95045
rect 21479 94981 21512 95045
rect 21304 94933 21512 94981
rect 788 90873 1322 90889
rect 788 90837 823 90873
rect 1279 90837 1322 90873
rect 788 90773 819 90837
rect 1283 90773 1322 90837
rect 788 90737 823 90773
rect 1279 90737 1322 90773
rect 788 90727 1322 90737
rect 1210 90653 36296 90665
rect 1210 90597 1805 90653
rect 1861 90597 1885 90653
rect 1941 90597 1965 90653
rect 2021 90597 2045 90653
rect 2101 90651 36296 90653
rect 2101 90597 24658 90651
rect 1210 90587 24658 90597
rect 24722 90587 24738 90651
rect 24802 90587 24818 90651
rect 24882 90587 24898 90651
rect 24962 90649 36296 90651
rect 24962 90587 34060 90649
rect 1210 90585 34060 90587
rect 34124 90585 34140 90649
rect 34204 90585 34220 90649
rect 34284 90585 34300 90649
rect 34364 90585 36296 90649
rect 1210 90571 36296 90585
rect 1206 90487 36296 90495
rect 1204 90482 36296 90487
rect 1204 90479 34594 90482
rect 1204 90474 27950 90479
rect 1204 90418 1455 90474
rect 1511 90418 1535 90474
rect 1591 90418 1615 90474
rect 1671 90423 27950 90474
rect 28006 90423 28030 90479
rect 28086 90423 34594 90479
rect 1671 90418 34594 90423
rect 34658 90418 34674 90482
rect 34738 90418 34754 90482
rect 34818 90418 34834 90482
rect 34898 90418 34914 90482
rect 34978 90418 34994 90482
rect 35058 90418 36296 90482
rect 1204 90401 36296 90418
rect 1204 90397 1502 90401
rect 1204 90331 2354 90333
rect 1200 90303 36296 90331
rect 1200 90287 35247 90303
rect 1200 89991 3053 90287
rect 3269 90286 35247 90287
rect 3269 90142 21333 90286
rect 21477 90142 35247 90286
rect 3269 89999 35247 90142
rect 35631 89999 36296 90303
rect 3269 89991 36296 89999
rect 1200 89931 36296 89991
rect 1210 89809 36296 89849
rect 1210 89539 2269 89809
rect 1224 89505 2269 89539
rect 2573 89801 36296 89809
rect 2573 89505 32676 89801
rect 1224 89497 32676 89505
rect 32820 89794 36296 89801
rect 32820 89497 35845 89794
rect 1224 89490 35845 89497
rect 36229 89490 36296 89794
rect 1224 89449 36296 89490
rect 0 87206 640 87223
rect 0 87070 51 87206
rect 587 87070 640 87206
rect 0 87021 640 87070
rect 33610 83515 34422 83571
rect 790 83267 1374 83298
rect 790 83123 843 83267
rect 1307 83123 1374 83267
rect 790 83100 1374 83123
rect 33610 83131 34064 83515
rect 34368 83131 34422 83515
rect 33610 83067 34422 83131
rect 0 82955 560 82961
rect 0 82953 1446 82955
rect 0 82933 1450 82953
rect 0 82789 854 82933
rect 1398 82789 1450 82933
rect 34580 82937 35070 82985
rect 0 82775 1450 82789
rect 806 82769 1450 82775
rect 21068 82856 21260 82905
rect 21068 82720 21099 82856
rect 21235 82720 21260 82856
rect 21068 81193 21260 82720
rect 34580 82633 34633 82937
rect 35017 82633 35070 82937
rect 34580 82577 35070 82633
rect 34798 82471 35212 82475
rect 36406 82471 36598 103383
rect 33004 82279 36598 82471
rect 34798 82277 35212 82279
rect 19202 77476 19814 77561
rect 19202 77020 19305 77476
rect 19681 77359 19814 77476
rect 21070 77359 21262 81092
rect 33630 80524 33806 80553
rect 33630 80300 33643 80524
rect 33787 80300 33806 80524
rect 33630 80288 33647 80300
rect 33783 80288 33806 80300
rect 33630 80257 33806 80288
rect 19681 77167 21262 77359
rect 19681 77020 19814 77167
rect 19202 76951 19814 77020
rect 23594 76575 24210 76587
rect 802 76571 33490 76575
rect 802 76542 33840 76571
rect 802 76398 854 76542
rect 1158 76519 33840 76542
rect 1158 76398 23659 76519
rect 802 76379 23659 76398
rect 806 76375 23659 76379
rect 23594 76063 23659 76375
rect 24115 76500 33840 76519
rect 24115 76436 33448 76500
rect 33512 76436 33528 76500
rect 33592 76436 33608 76500
rect 33672 76436 33688 76500
rect 33752 76436 33768 76500
rect 33832 76436 33840 76500
rect 24115 76375 33840 76436
rect 24115 76063 24210 76375
rect 33410 76361 33840 76375
rect 32200 76233 32752 76235
rect 23594 75993 24210 76063
rect 32198 76144 32762 76233
rect 0 75873 1624 75883
rect 32198 75873 32252 76144
rect 0 75768 32252 75873
rect 32708 75768 32762 76144
rect 0 75695 32762 75768
rect 0 75681 32752 75695
rect 32200 75677 32752 75681
rect 34048 75471 34374 75491
rect 34048 75007 34059 75471
rect 34363 75007 34374 75471
rect 34048 74987 34374 75007
rect 34598 74688 35030 74689
rect 34598 74224 34622 74688
rect 35006 74224 35030 74688
rect 34598 74223 35030 74224
rect 35258 73866 35664 73871
rect 35258 73402 35269 73866
rect 35653 73402 35664 73866
rect 35258 73397 35664 73402
rect 35826 73063 36246 73091
rect 35826 72599 35844 73063
rect 36228 72599 36246 73063
rect 35826 72571 36246 72599
rect 0 64171 2356 64347
rect 0 57445 2360 57621
rect 0 50729 2352 50905
rect 0 44035 2364 44211
rect 0 37265 2368 37441
rect 0 36353 2356 36529
rect 0 35887 2346 36063
rect 0 30279 2356 30455
rect 0 23573 2364 23749
rect 0 16853 2360 17029
rect 0 10151 2352 10327
rect 0 3373 2356 3549
rect 0 2230 888 2235
rect 1212 2230 2650 2231
rect 0 1835 2650 2230
rect 1212 1833 2650 1835
rect 0 1697 888 1699
rect 0 1299 2644 1697
rect 0 1195 924 1199
rect 0 807 2688 1195
rect 0 255 2686 635
<< via3 >>
rect 27895 99499 28119 99503
rect 27895 99043 27899 99499
rect 27899 99043 28115 99499
rect 28115 99043 28119 99499
rect 27895 99039 28119 99043
rect 21335 94981 21399 95045
rect 21415 94981 21479 95045
rect 819 90773 823 90837
rect 823 90773 883 90837
rect 899 90773 963 90837
rect 979 90773 1043 90837
rect 1059 90773 1123 90837
rect 1139 90773 1203 90837
rect 1219 90773 1279 90837
rect 1279 90773 1283 90837
rect 24658 90587 24722 90651
rect 24738 90587 24802 90651
rect 24818 90587 24882 90651
rect 24898 90587 24962 90651
rect 34060 90585 34124 90649
rect 34140 90585 34204 90649
rect 34220 90585 34284 90649
rect 34300 90585 34364 90649
rect 34594 90418 34658 90482
rect 34674 90418 34738 90482
rect 34754 90418 34818 90482
rect 34834 90418 34898 90482
rect 34914 90418 34978 90482
rect 34994 90418 35058 90482
rect 21333 90142 21477 90286
rect 35247 89999 35631 90303
rect 2269 89505 2573 89809
rect 32676 89497 32820 89801
rect 35845 89490 36229 89794
rect 843 83263 1307 83267
rect 843 83127 847 83263
rect 847 83127 1303 83263
rect 1303 83127 1307 83263
rect 843 83123 1307 83127
rect 34064 83131 34368 83515
rect 854 82929 1398 82933
rect 854 82793 858 82929
rect 858 82793 1394 82929
rect 1394 82793 1398 82929
rect 854 82789 1398 82793
rect 34633 82933 35017 82937
rect 34633 82637 34637 82933
rect 34637 82637 35013 82933
rect 35013 82637 35017 82933
rect 34633 82633 35017 82637
rect 33643 80424 33787 80524
rect 33643 80300 33647 80424
rect 33647 80300 33783 80424
rect 33783 80300 33787 80424
rect 854 76398 1158 76542
rect 33448 76436 33512 76500
rect 33528 76436 33592 76500
rect 33608 76436 33672 76500
rect 33688 76436 33752 76500
rect 33768 76436 33832 76500
rect 34059 75007 34363 75471
rect 34622 74224 35006 74688
rect 35269 73402 35653 73866
rect 35844 72599 36228 73063
<< metal4 >>
rect 27894 99503 28120 99537
rect 27894 99039 27895 99503
rect 28119 99039 28120 99503
rect 27894 99005 28120 99039
rect 21304 95045 21512 95085
rect 21304 94981 21335 95045
rect 21399 94981 21415 95045
rect 21479 94981 21512 95045
rect 21304 94933 21512 94981
rect 788 90837 1322 90889
rect 788 90773 819 90837
rect 883 90773 899 90837
rect 963 90773 979 90837
rect 1043 90773 1059 90837
rect 1123 90773 1139 90837
rect 1203 90773 1219 90837
rect 1283 90773 1322 90837
rect 788 90727 1322 90773
rect 792 84058 992 90727
rect 21304 90286 21510 94933
rect 24650 90651 24970 98747
rect 24650 90587 24658 90651
rect 24722 90587 24738 90651
rect 24802 90587 24818 90651
rect 24882 90587 24898 90651
rect 24962 90587 24970 90651
rect 24650 90573 24970 90587
rect 34016 90649 34412 90663
rect 34016 90585 34060 90649
rect 34124 90585 34140 90649
rect 34204 90585 34220 90649
rect 34284 90585 34300 90649
rect 34364 90585 34412 90649
rect 21304 90142 21333 90286
rect 21477 90142 21510 90286
rect 2202 89809 2626 89849
rect 2202 89505 2269 89809
rect 2573 89505 2626 89809
rect 2202 89154 2626 89505
rect 2202 88881 2628 89154
rect 2208 88524 2628 88881
rect 21304 87952 21510 90142
rect 32627 89801 32861 89848
rect 32627 89497 32676 89801
rect 32820 89497 32861 89801
rect 32627 87932 32861 89497
rect 776 83632 992 84058
rect 792 83298 992 83632
rect 34016 83587 34412 90585
rect 34588 90482 35066 90672
rect 34588 90418 34594 90482
rect 34658 90418 34674 90482
rect 34738 90418 34754 90482
rect 34818 90418 34834 90482
rect 34898 90418 34914 90482
rect 34978 90418 34994 90482
rect 35058 90418 35066 90482
rect 34016 83515 34428 83587
rect 790 83267 1374 83298
rect 790 83123 843 83267
rect 1307 83123 1374 83267
rect 790 83100 1374 83123
rect 34016 83131 34064 83515
rect 34368 83131 34428 83515
rect 792 83098 1372 83100
rect 792 83096 992 83098
rect 34016 83055 34428 83131
rect 804 82953 1012 82959
rect 804 82933 1450 82953
rect 804 82789 854 82933
rect 1398 82789 1450 82933
rect 804 82769 1450 82789
rect 804 76575 1012 82769
rect 33630 80524 33810 80555
rect 33630 80300 33643 80524
rect 33787 80300 33810 80524
rect 33630 80257 33810 80300
rect 802 76542 1216 76575
rect 33630 76571 33808 80257
rect 802 76398 854 76542
rect 1158 76398 1216 76542
rect 802 76379 1216 76398
rect 33410 76500 33840 76571
rect 33410 76436 33448 76500
rect 33512 76436 33528 76500
rect 33592 76436 33608 76500
rect 33672 76436 33688 76500
rect 33752 76436 33768 76500
rect 33832 76436 33840 76500
rect 33410 76361 33840 76436
rect 34016 75471 34412 83055
rect 34016 75007 34059 75471
rect 34363 75007 34412 75471
rect 34016 74921 34412 75007
rect 34588 82989 35066 90418
rect 35204 90303 35682 90664
rect 35204 89999 35247 90303
rect 35631 89999 35682 90303
rect 34588 82937 35070 82989
rect 34588 82633 34633 82937
rect 35017 82633 35070 82937
rect 34588 82577 35070 82633
rect 34588 74688 35066 82577
rect 34588 74224 34622 74688
rect 35006 74224 35066 74688
rect 34588 74150 35066 74224
rect 35204 73866 35682 89999
rect 35204 73402 35269 73866
rect 35653 73402 35682 73866
rect 35204 73352 35682 73402
rect 35806 89794 36284 90667
rect 35806 89490 35845 89794
rect 36229 89490 36284 89794
rect 35806 73063 36284 89490
rect 35806 72599 35844 73063
rect 36228 72599 36284 73063
rect 35806 72550 36284 72599
use EF_AMUX0801WISO  EF_AMUX0801WISO_0
timestamp 1699520070
transform 1 0 1516 0 -1 101767
box -306 -2006 33704 11044
use EF_DACSCA1001  EF_DACSCA1001_0
timestamp 1699520070
transform 1 0 2156 0 1 7338
box -946 -7090 66618 68998
use EF_R2RVCE  EF_R2RVCE_0
timestamp 1699520070
transform 1 0 21872 0 1 78162
box -804 -1465 11921 11144
use sample_and_hold  sample_and_hold_0
timestamp 1699520070
transform 1 0 1174 0 1 78112
box 0 -114 19469 11183
<< labels >>
flabel metal1 s 1174 87018 1374 87218 0 FreeSans 30 0 0 0 HOLD
port 1 nsew
flabel metal2 s 27962 103465 28050 103773 0 FreeSans 150 0 0 0 VIN[0]
port 2 nsew
flabel metal2 s 24516 103467 24612 103773 0 FreeSans 150 0 0 0 VIN[1]
port 3 nsew
flabel metal2 s 21214 103467 21310 103773 0 FreeSans 150 0 0 0 VIN[2]
port 4 nsew
flabel metal2 s 17840 103467 17936 103773 0 FreeSans 150 0 0 0 VIN[3]
port 5 nsew
flabel metal2 s 14528 103465 14618 103773 0 FreeSans 150 0 0 0 VIN[4]
port 6 nsew
flabel metal2 s 11230 103465 11320 103773 0 FreeSans 150 0 0 0 VIN[5]
port 7 nsew
flabel metal2 s 7828 103473 7918 103773 0 FreeSans 150 0 0 0 VIN[6]
port 8 nsew
flabel metal2 s 4424 103475 4520 103773 0 FreeSans 150 0 0 0 VIN[7]
port 9 nsew
flabel metal3 s 0 87021 640 87223 0 FreeSans 600 0 0 0 HOLD
port 1 nsew
flabel metal3 s 0 82775 560 82961 0 FreeSans 600 0 0 0 EN
port 10 nsew
flabel metal3 s 0 75681 500 75883 0 FreeSans 600 0 0 0 RST
port 11 nsew
flabel metal3 s 0 64171 554 64347 0 FreeSans 600 0 0 0 DATA[9]
port 12 nsew
flabel metal3 s 0 57445 648 57621 0 FreeSans 600 0 0 0 DATA[8]
port 13 nsew
flabel metal3 s 0 50729 648 50905 0 FreeSans 600 0 0 0 DATA[7]
port 14 nsew
flabel metal3 s 0 44035 648 44211 0 FreeSans 600 0 0 0 DATA[6]
port 15 nsew
flabel metal3 s 0 37265 648 37441 0 FreeSans 600 0 0 0 DATA[5]
port 16 nsew
flabel metal3 s 0 30279 648 30455 0 FreeSans 600 0 0 0 DATA[0]
port 17 nsew
flabel metal3 s 0 23573 648 23749 0 FreeSans 600 0 0 0 DATA[1]
port 18 nsew
flabel metal3 s 0 16853 648 17029 0 FreeSans 600 0 0 0 DATA[2]
port 19 nsew
flabel metal3 s 0 10151 648 10327 0 FreeSans 600 0 0 0 DATA[3]
port 20 nsew
flabel metal3 s 0 3373 648 3549 0 FreeSans 600 0 0 0 DATA[4]
port 21 nsew
flabel metal3 s 0 1299 888 1699 0 FreeSans 600 0 0 0 DVSS
port 22 nsew
flabel metal3 s 0 1835 888 2235 0 FreeSans 600 0 0 0 DVDD
port 23 nsew
flabel metal3 s 0 807 924 1199 0 FreeSans 600 0 0 0 VDD
port 24 nsew
flabel metal3 s 0 255 940 635 0 FreeSans 600 0 0 0 VSS
port 25 nsew
flabel metal3 s 0 36353 658 36529 0 FreeSans 600 0 0 0 VH
port 26 nsew
flabel metal3 s 0 35887 658 36063 0 FreeSans 600 0 0 0 VL
port 27 nsew
flabel metal2 s 35196 103589 35256 103773 0 FreeSans 600 0 0 0 B[0]
port 28 nsew
flabel metal2 s 35342 103585 35402 103773 0 FreeSans 600 0 0 0 B[1]
port 29 nsew
flabel metal2 s 35488 103585 35548 103773 0 FreeSans 600 0 0 0 B[2]
port 30 nsew
flabel metal2 s 36404 103333 36598 103773 0 FreeSans 600 0 0 0 CMP
port 31 nsew
<< end >>
