magic
tech sky130A
magscale 1 2
timestamp 1694031861
<< metal1 >>
rect 3400 7042 27400 7264
rect 5846 3328 6036 4158
rect 9298 3336 9488 4166
rect 12636 3274 12826 4104
rect 16062 3314 16252 4144
rect 19450 3296 19640 4126
rect 22880 3306 23070 4136
rect 26236 3336 26426 4166
rect 29674 3328 29878 4184
rect 30208 3444 30676 3454
rect 30208 3407 30690 3444
rect 30208 2971 30271 3407
rect 30579 2971 30690 3407
rect 30208 2902 30690 2971
rect 13810 1499 14024 1508
rect 7020 1481 7234 1492
rect 3604 1466 3818 1478
rect 3604 1286 3612 1466
rect 3792 1286 3818 1466
rect 7020 1301 7035 1481
rect 7215 1301 7234 1481
rect 7020 1286 7234 1301
rect 10400 1488 10614 1496
rect 10400 1308 10413 1488
rect 10593 1308 10614 1488
rect 10400 1290 10614 1308
rect 13810 1319 13856 1499
rect 13972 1319 14024 1499
rect 20616 1498 20850 1504
rect 13810 1302 14024 1319
rect 17194 1484 17408 1486
rect 17194 1480 17416 1484
rect 17194 1300 17219 1480
rect 17399 1300 17416 1480
rect 20616 1318 20642 1498
rect 20822 1318 20850 1498
rect 27412 1494 27626 1504
rect 20616 1302 20850 1318
rect 23994 1479 24208 1486
rect 17194 1296 17416 1300
rect 3604 1272 3818 1286
rect 17194 1280 17408 1296
rect 20622 1290 20836 1302
rect 23994 1299 24014 1479
rect 24194 1299 24208 1479
rect 23994 1280 24208 1299
rect 27412 1314 27431 1494
rect 27611 1314 27626 1494
rect 27412 1298 27626 1314
rect 30212 1186 30690 2902
rect 30058 1154 30690 1186
rect 6246 966 30690 1154
rect 30058 962 30690 966
rect 30058 952 30638 962
<< via1 >>
rect 30271 2971 30579 3407
rect 3612 1286 3792 1466
rect 7035 1301 7215 1481
rect 10413 1308 10593 1488
rect 13856 1319 13972 1499
rect 17219 1300 17399 1480
rect 20642 1318 20822 1498
rect 24014 1299 24194 1479
rect 27431 1314 27611 1494
<< metal2 >>
rect 30208 3417 30676 3454
rect 30208 3407 30277 3417
rect 30573 3407 30676 3417
rect 30208 2971 30271 3407
rect 30579 2971 30676 3407
rect 30208 2961 30277 2971
rect 30573 2961 30676 2971
rect 30208 2902 30676 2961
rect 13796 1499 14026 1516
rect 6998 1481 7260 1496
rect 3594 1466 3810 1474
rect 3594 1286 3612 1466
rect 3792 1286 3810 1466
rect 3594 -1500 3810 1286
rect 6998 1301 7035 1481
rect 7215 1301 7260 1481
rect 6998 -1188 7260 1301
rect 10396 1488 10616 1498
rect 10396 1308 10413 1488
rect 10593 1308 10616 1488
rect 10396 -900 10616 1308
rect 13796 1319 13856 1499
rect 13972 1319 14026 1499
rect 20600 1504 20848 1510
rect 20600 1498 20850 1504
rect 13796 -590 14026 1319
rect 17196 1480 17420 1490
rect 17196 1300 17219 1480
rect 17399 1300 17420 1480
rect 17196 -278 17420 1300
rect 20600 1318 20642 1498
rect 20822 1318 20850 1498
rect 23998 1490 24214 1496
rect 27406 1494 27624 1508
rect 20600 1302 20850 1318
rect 23992 1479 24220 1490
rect 20600 8 20848 1302
rect 23992 1299 24014 1479
rect 24194 1299 24220 1479
rect 23992 1290 24220 1299
rect 27406 1314 27431 1494
rect 27611 1314 27624 1494
rect 23998 718 24214 1290
rect 23994 620 24214 718
rect 27406 630 27624 1314
rect 23994 304 24212 620
rect 27400 584 27828 630
rect 27400 448 27464 584
rect 27760 448 27828 584
rect 27400 400 27828 448
rect 27406 391 27624 400
rect 23994 302 24440 304
rect 23984 285 24454 302
rect 23984 149 24024 285
rect 24400 149 24454 285
rect 23984 126 24454 149
rect 23994 112 24440 126
rect 23994 108 24212 112
rect 20600 -26 20992 8
rect 20600 -162 20647 -26
rect 20943 -162 20992 -26
rect 20600 -196 20992 -162
rect 17196 -316 17624 -278
rect 17196 -452 17226 -316
rect 17602 -452 17624 -316
rect 17196 -488 17624 -452
rect 13796 -622 14258 -590
rect 13796 -758 13836 -622
rect 14212 -758 14258 -622
rect 13796 -790 14258 -758
rect 13796 -791 14026 -790
rect 10382 -926 10812 -900
rect 10382 -1062 10404 -926
rect 10780 -1062 10812 -926
rect 10382 -1096 10812 -1062
rect 6998 -1231 7512 -1188
rect 6998 -1367 7074 -1231
rect 7450 -1367 7512 -1231
rect 6998 -1405 7512 -1367
rect 7000 -1406 7512 -1405
rect 3594 -1533 4104 -1500
rect 3594 -1669 3670 -1533
rect 4046 -1669 4104 -1533
rect 3594 -1712 4104 -1669
rect 3594 -1716 3810 -1712
<< via2 >>
rect 30277 3407 30573 3417
rect 30277 2971 30573 3407
rect 30277 2961 30573 2971
rect 27464 448 27760 584
rect 24024 149 24400 285
rect 20647 -162 20943 -26
rect 17226 -452 17602 -316
rect 13836 -758 14212 -622
rect 10404 -1062 10780 -926
rect 7074 -1367 7450 -1231
rect 3670 -1669 4046 -1533
<< metal3 >>
rect 6326 4812 26916 5056
rect 31594 4562 31656 4752
rect 34178 4566 34240 4720
rect 36898 4594 36962 4776
rect 26744 4016 27012 4074
rect 26744 3632 26808 4016
rect 26952 3632 27012 4016
rect 26744 1697 27012 3632
rect 30208 3421 30676 3454
rect 30208 2957 30273 3421
rect 30577 2957 30676 3421
rect 30208 2902 30676 2957
rect 6461 1539 27012 1697
rect 26744 1536 27012 1539
rect 30778 644 30838 816
rect 27400 588 27828 630
rect 27400 444 27460 588
rect 27764 444 27828 588
rect 27400 400 27828 444
rect 30388 586 30872 644
rect 30388 442 30440 586
rect 30824 442 30872 586
rect 30388 392 30872 442
rect 31600 552 31900 704
rect 23996 302 24440 304
rect 23984 289 24454 302
rect 23984 145 24020 289
rect 24404 145 24454 289
rect 23984 126 24454 145
rect 31600 282 31902 552
rect 31600 138 31638 282
rect 31862 138 31902 282
rect 23996 112 24440 126
rect 31600 112 31902 138
rect 20600 -22 20992 8
rect 20600 -166 20643 -22
rect 20947 -166 20992 -22
rect 20600 -196 20992 -166
rect 32540 -26 32840 696
rect 33774 672 33832 678
rect 33768 670 33832 672
rect 32540 -170 32580 -26
rect 32804 -170 32840 -26
rect 32540 -196 32840 -170
rect 33642 -58 33930 670
rect 33642 -274 33936 -58
rect 17200 -312 17624 -278
rect 17200 -456 17222 -312
rect 17606 -456 17624 -312
rect 17200 -488 17624 -456
rect 33636 -310 33936 -274
rect 33636 -454 33677 -310
rect 33901 -454 33936 -310
rect 33636 -486 33936 -454
rect 13796 -618 14258 -590
rect 13796 -762 13832 -618
rect 14216 -762 14258 -618
rect 13796 -790 14258 -762
rect 34620 -619 34892 708
rect 37514 694 37578 708
rect 34620 -763 34645 -619
rect 34869 -763 34892 -619
rect 34620 -786 34892 -763
rect 10382 -922 10812 -900
rect 10382 -1066 10400 -922
rect 10784 -1066 10812 -922
rect 10382 -1096 10812 -1066
rect 35602 -916 35886 690
rect 36684 574 36974 678
rect 36684 280 36986 574
rect 35602 -1060 35632 -916
rect 35856 -1060 35886 -916
rect 35602 -1082 35886 -1060
rect 7000 -1227 7512 -1188
rect 7000 -1371 7070 -1227
rect 7454 -1371 7512 -1227
rect 7000 -1406 7512 -1371
rect 36694 -1228 36986 280
rect 36694 -1372 36742 -1228
rect 36966 -1372 36986 -1228
rect 36694 -1410 36986 -1372
rect 3610 -1529 4104 -1500
rect 3610 -1673 3666 -1529
rect 4050 -1673 4104 -1529
rect 3610 -1712 4104 -1673
rect 37410 -1530 37670 694
rect 37410 -1674 37470 -1530
rect 37614 -1674 37670 -1530
rect 37410 -1700 37670 -1674
<< via3 >>
rect 26808 3632 26952 4016
rect 30273 3417 30577 3421
rect 30273 2961 30277 3417
rect 30277 2961 30573 3417
rect 30573 2961 30577 3417
rect 30273 2957 30577 2961
rect 27460 584 27764 588
rect 27460 448 27464 584
rect 27464 448 27760 584
rect 27760 448 27764 584
rect 27460 444 27764 448
rect 30440 442 30824 586
rect 24020 285 24404 289
rect 24020 149 24024 285
rect 24024 149 24400 285
rect 24400 149 24404 285
rect 24020 145 24404 149
rect 31638 138 31862 282
rect 20643 -26 20947 -22
rect 20643 -162 20647 -26
rect 20647 -162 20943 -26
rect 20943 -162 20947 -26
rect 20643 -166 20947 -162
rect 32580 -170 32804 -26
rect 17222 -316 17606 -312
rect 17222 -452 17226 -316
rect 17226 -452 17602 -316
rect 17602 -452 17606 -316
rect 17222 -456 17606 -452
rect 33677 -454 33901 -310
rect 13832 -622 14216 -618
rect 13832 -758 13836 -622
rect 13836 -758 14212 -622
rect 14212 -758 14216 -622
rect 13832 -762 14216 -758
rect 34645 -763 34869 -619
rect 10400 -926 10784 -922
rect 10400 -1062 10404 -926
rect 10404 -1062 10780 -926
rect 10780 -1062 10784 -926
rect 10400 -1066 10784 -1062
rect 35632 -1060 35856 -916
rect 7070 -1231 7454 -1227
rect 7070 -1367 7074 -1231
rect 7074 -1367 7450 -1231
rect 7450 -1367 7454 -1231
rect 7070 -1371 7454 -1367
rect 36742 -1372 36966 -1228
rect 3666 -1533 4050 -1529
rect 3666 -1669 3670 -1533
rect 3670 -1669 4046 -1533
rect 4046 -1669 4050 -1533
rect 3666 -1673 4050 -1669
rect 37470 -1674 37614 -1530
<< metal4 >>
rect 26748 4074 27000 4078
rect 27082 4074 31110 4080
rect 26744 4016 31110 4074
rect 26744 3760 26808 4016
rect 26748 3632 26808 3760
rect 26952 3760 31110 4016
rect 26952 3632 27000 3760
rect 26748 3574 27000 3632
rect 30208 3444 30676 3454
rect 30208 3421 31050 3444
rect 30208 2957 30273 3421
rect 30577 3126 31050 3421
rect 30577 2957 30676 3126
rect 30208 2902 30676 2957
rect 30388 636 30872 644
rect 27378 588 30872 636
rect 27378 444 27460 588
rect 27764 586 30872 588
rect 27764 444 30440 586
rect 27378 442 30440 444
rect 30824 442 30872 586
rect 27378 392 30872 442
rect 31600 304 31900 308
rect 23992 302 31900 304
rect 23984 289 31900 302
rect 23984 145 24020 289
rect 24404 282 31900 289
rect 24404 145 31638 282
rect 23984 138 31638 145
rect 31862 138 31900 282
rect 23984 126 31900 138
rect 23992 114 31900 126
rect 31600 112 31900 114
rect 20602 -22 32842 8
rect 20602 -166 20643 -22
rect 20947 -26 32842 -22
rect 20947 -166 32580 -26
rect 20602 -170 32580 -166
rect 32804 -170 32842 -26
rect 20602 -198 32842 -170
rect 17186 -310 33960 -282
rect 17186 -312 33677 -310
rect 17186 -456 17222 -312
rect 17606 -454 33677 -312
rect 33901 -454 33960 -310
rect 17606 -456 33960 -454
rect 17186 -490 33960 -456
rect 13694 -618 34912 -592
rect 13694 -762 13832 -618
rect 14216 -619 34912 -618
rect 14216 -762 34645 -619
rect 13694 -763 34645 -762
rect 34869 -763 34912 -619
rect 13694 -790 34912 -763
rect 10394 -916 35888 -906
rect 10394 -922 35632 -916
rect 10394 -1066 10400 -922
rect 10784 -1060 35632 -922
rect 35856 -1060 35888 -916
rect 10784 -1066 35888 -1060
rect 10394 -1096 35888 -1066
rect 6992 -1227 36990 -1204
rect 6992 -1371 7070 -1227
rect 7454 -1228 36990 -1227
rect 7454 -1371 36742 -1228
rect 6992 -1372 36742 -1371
rect 36966 -1372 36990 -1228
rect 6992 -1410 36990 -1372
rect 3548 -1529 37700 -1504
rect 3548 -1673 3666 -1529
rect 4050 -1530 37700 -1529
rect 4050 -1673 37470 -1530
rect 3548 -1674 37470 -1673
rect 37614 -1674 37700 -1530
rect 3548 -1710 37700 -1674
use array_2ls_2tgm  array_2ls_2tgm_0
timestamp 1694031861
transform 1 0 30200 0 1 614
box -6569 341 -73 6588
use array_2ls_2tgm  array_2ls_2tgm_1
timestamp 1694031861
transform 1 0 9814 0 1 602
box -6569 341 -73 6588
use array_2ls_2tgm  array_2ls_2tgm_2
timestamp 1694031861
transform 1 0 16598 0 1 620
box -6569 341 -73 6588
use array_2ls_2tgm  array_2ls_2tgm_3
timestamp 1694031861
transform 1 0 23406 0 1 614
box -6569 341 -73 6588
use decoder3to8  decoder3to8_0
timestamp 1694031861
transform 0 1 30335 -1 0 4644
box -222 426 4178 7249
<< labels >>
flabel metal3 s 36912 4658 36938 4706 0 FreeSans 244 0 0 0 B[0]
port 1 nsew
flabel metal3 s 34194 4628 34224 4694 0 FreeSans 244 0 0 0 B[1]
port 2 nsew
flabel metal3 s 31608 4622 31638 4678 0 FreeSans 244 0 0 0 B[2]
port 3 nsew
flabel metal1 s 29726 3630 29782 3680 0 FreeSans 244 0 0 0 VIN[0]
port 4 nsew
flabel metal1 s 26288 3812 26350 3888 0 FreeSans 244 0 0 0 VIN[1]
port 5 nsew
flabel metal1 s 22926 3674 22990 3732 0 FreeSans 244 0 0 0 VIN[2]
port 6 nsew
flabel metal1 s 19532 3790 19590 3872 0 FreeSans 244 0 0 0 VIN[3]
port 7 nsew
flabel metal1 s 16138 3730 16206 3796 0 FreeSans 244 0 0 0 VIN[4]
port 8 nsew
flabel metal1 s 12700 3668 12754 3760 0 FreeSans 244 0 0 0 VIN[5]
port 9 nsew
flabel metal1 s 9350 3712 9414 3750 0 FreeSans 244 0 0 0 VIN[6]
port 10 nsew
flabel metal1 s 5904 3630 5980 3710 0 FreeSans 244 0 0 0 VIN[7]
port 11 nsew
flabel metal1 s 29856 1044 29902 1098 0 FreeSans 244 0 0 0 VSS
port 12 nsew
flabel metal1 s 23200 7078 23258 7160 0 FreeSans 244 0 0 0 VO
port 13 nsew
flabel metal3 s 12806 4864 12866 4970 0 FreeSans 244 0 0 0 VDD3V3
port 14 nsew
flabel metal3 s 23384 1578 23460 1646 0 FreeSans 244 0 0 0 VDD1V8
port 15 nsew
<< end >>
