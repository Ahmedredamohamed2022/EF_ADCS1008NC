VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO EF_ADCS1008NC
  CLASS BLOCK ;
  FOREIGN EF_ADCS1008NC ;
  ORIGIN 15.140 4.960 ;
  SIZE 178.485 BY 487.030 ;
  PIN DVSS
    ANTENNAGATEAREA 74.759102 ;
    ANTENNADIFFAREA 816.096802 ;
    PORT
      LAYER met3 ;
        RECT 5.400 -1.830 6.090 -1.550 ;
    END
  END DVSS
  PIN DVDD
    ANTENNAGATEAREA 47.261497 ;
    ANTENNADIFFAREA 92.613647 ;
    PORT
      LAYER met3 ;
        RECT 4.430 0.430 5.120 1.140 ;
    END
  END DVDD
  PIN VDD
    ANTENNAGATEAREA 100.000000 ;
    ANTENNADIFFAREA 2017.665894 ;
    PORT
      LAYER met3 ;
        RECT 4.100 -4.300 4.790 -3.590 ;
    END
  END VDD
  PIN VH
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met3 ;
        RECT 3.030 29.620 3.460 30.540 ;
    END
  END VH
  PIN VL
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met3 ;
        RECT 1.250 31.130 1.560 32.020 ;
    END
  END VL
  PIN VSS
    ANTENNAGATEAREA 130.000000 ;
    ANTENNADIFFAREA 530.402893 ;
    PORT
      LAYER met3 ;
        RECT 96.070 346.940 97.480 348.330 ;
    END
  END VSS
  PIN EN
    ANTENNAGATEAREA 1.500000 ;
    ANTENNADIFFAREA 1.080000 ;
    PORT
      LAYER met1 ;
        RECT 92.350 284.450 92.650 284.820 ;
    END
  END EN
  PIN RST
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER met3 ;
        RECT 127.770 316.630 128.510 317.080 ;
    END
  END RST
  PIN HOLD
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT -2.890 405.500 -2.620 405.800 ;
    END
  END HOLD
  PIN CMP
    ANTENNADIFFAREA 0.492900 ;
    PORT
      LAYER met2 ;
        RECT 129.380 422.350 130.660 423.270 ;
    END
  END CMP
  PIN DATA[0]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met1 ;
        RECT 5.770 13.720 6.190 14.660 ;
    END
  END DATA[0]
  PIN DATA[1]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met1 ;
        RECT 5.770 49.740 6.070 50.480 ;
    END
  END DATA[1]
  PIN DATA[2]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met1 ;
        RECT 5.790 83.250 6.190 84.160 ;
    END
  END DATA[2]
  PIN DATA[3]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met1 ;
        RECT 5.790 117.860 6.200 118.700 ;
    END
  END DATA[3]
  PIN DATA[4]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met1 ;
        RECT 5.970 152.860 6.270 153.910 ;
    END
  END DATA[4]
  PIN DATA[5]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met1 ;
        RECT 5.790 184.510 6.150 185.350 ;
    END
  END DATA[5]
  PIN DATA[6]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met1 ;
        RECT 5.670 219.460 6.050 220.550 ;
    END
  END DATA[6]
  PIN DATA[7]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met1 ;
        RECT 5.740 252.410 6.200 253.470 ;
    END
  END DATA[7]
  PIN DATA[8]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met1 ;
        RECT 5.940 285.500 6.270 286.030 ;
    END
  END DATA[8]
  PIN DATA[9]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met1 ;
        RECT 5.940 321.970 6.250 322.790 ;
    END
  END DATA[9]
  PIN B[0]
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 159.380 449.530 159.610 449.700 ;
    END
  END B[0]
  PIN B[1]
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 145.870 449.620 146.050 449.800 ;
    END
  END B[1]
  PIN B[2]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 132.890 449.450 133.010 449.540 ;
    END
  END B[2]
  PIN VIN[7]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met1 ;
        RECT 4.450 456.730 4.840 457.170 ;
    END
  END VIN[7]
  PIN VIN[6]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met1 ;
        RECT 21.650 457.250 21.870 457.660 ;
    END
  END VIN[6]
  PIN VIN[5]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met1 ;
        RECT 38.450 457.220 38.610 457.370 ;
    END
  END VIN[5]
  PIN VIN[4]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met1 ;
        RECT 55.430 457.520 55.760 458.070 ;
    END
  END VIN[4]
  PIN VIN[3]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met1 ;
        RECT 72.320 457.170 72.690 457.400 ;
    END
  END VIN[3]
  PIN VIN[2]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met1 ;
        RECT 89.640 457.510 89.980 457.790 ;
    END
  END VIN[2]
  PIN VIN[1]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met1 ;
        RECT 106.240 457.110 106.700 457.250 ;
    END
  END VIN[1]
  PIN VIN[0]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met1 ;
        RECT 123.650 457.490 123.790 457.790 ;
    END
  END VIN[0]
  OBS
      LAYER li1 ;
        RECT -8.600 7.615 161.965 469.590 ;
      LAYER met1 ;
        RECT -15.090 458.350 162.120 469.590 ;
        RECT -15.090 457.940 55.150 458.350 ;
        RECT -15.090 457.450 21.370 457.940 ;
        RECT -15.090 456.450 4.170 457.450 ;
        RECT 5.120 456.970 21.370 457.450 ;
        RECT 22.150 457.650 55.150 457.940 ;
        RECT 22.150 456.970 38.170 457.650 ;
        RECT 5.120 456.940 38.170 456.970 ;
        RECT 38.890 457.240 55.150 457.650 ;
        RECT 56.040 458.070 162.120 458.350 ;
        RECT 56.040 457.680 89.360 458.070 ;
        RECT 56.040 457.240 72.040 457.680 ;
        RECT 38.890 456.940 72.040 457.240 ;
        RECT 5.120 456.890 72.040 456.940 ;
        RECT 72.970 457.230 89.360 457.680 ;
        RECT 90.260 457.530 123.370 458.070 ;
        RECT 90.260 457.230 105.960 457.530 ;
        RECT 72.970 456.890 105.960 457.230 ;
        RECT 5.120 456.830 105.960 456.890 ;
        RECT 106.980 457.210 123.370 457.530 ;
        RECT 124.070 457.210 162.120 458.070 ;
        RECT 106.980 456.830 162.120 457.210 ;
        RECT 5.120 456.450 162.120 456.830 ;
        RECT -15.090 406.080 162.120 456.450 ;
        RECT -15.090 405.220 -3.170 406.080 ;
        RECT -2.340 405.220 162.120 406.080 ;
        RECT -15.090 323.070 162.120 405.220 ;
        RECT -15.090 321.690 5.660 323.070 ;
        RECT 6.530 321.690 162.120 323.070 ;
        RECT -15.090 286.310 162.120 321.690 ;
        RECT -15.090 285.220 5.660 286.310 ;
        RECT 6.550 285.220 162.120 286.310 ;
        RECT -15.090 285.100 162.120 285.220 ;
        RECT -15.090 284.170 92.070 285.100 ;
        RECT 92.930 284.170 162.120 285.100 ;
        RECT -15.090 253.750 162.120 284.170 ;
        RECT -15.090 252.130 5.460 253.750 ;
        RECT 6.480 252.130 162.120 253.750 ;
        RECT -15.090 220.830 162.120 252.130 ;
        RECT -15.090 219.180 5.390 220.830 ;
        RECT 6.330 219.180 162.120 220.830 ;
        RECT -15.090 185.630 162.120 219.180 ;
        RECT -15.090 184.230 5.510 185.630 ;
        RECT 6.430 184.230 162.120 185.630 ;
        RECT -15.090 154.190 162.120 184.230 ;
        RECT -15.090 152.580 5.690 154.190 ;
        RECT 6.550 152.580 162.120 154.190 ;
        RECT -15.090 118.980 162.120 152.580 ;
        RECT -15.090 117.580 5.510 118.980 ;
        RECT 6.480 117.580 162.120 118.980 ;
        RECT -15.090 84.440 162.120 117.580 ;
        RECT -15.090 82.970 5.510 84.440 ;
        RECT 6.470 82.970 162.120 84.440 ;
        RECT -15.090 50.760 162.120 82.970 ;
        RECT -15.090 49.460 5.490 50.760 ;
        RECT 6.350 49.460 162.120 50.760 ;
        RECT -15.090 14.940 162.120 49.460 ;
        RECT -15.090 13.440 5.490 14.940 ;
        RECT 6.470 13.440 162.120 14.940 ;
        RECT -15.090 5.090 162.120 13.440 ;
      LAYER met2 ;
        RECT -15.100 423.550 162.765 482.070 ;
        RECT -15.100 422.070 129.100 423.550 ;
        RECT 130.940 422.070 162.765 423.550 ;
        RECT -15.100 3.010 162.765 422.070 ;
      LAYER met3 ;
        RECT -15.140 450.200 163.195 482.050 ;
        RECT -15.140 449.940 145.470 450.200 ;
        RECT -15.140 449.050 132.490 449.940 ;
        RECT 133.410 449.220 145.470 449.940 ;
        RECT 146.450 450.100 163.195 450.200 ;
        RECT 146.450 449.220 158.980 450.100 ;
        RECT 133.410 449.130 158.980 449.220 ;
        RECT 160.010 449.130 163.195 450.100 ;
        RECT 133.410 449.050 163.195 449.130 ;
        RECT -15.140 348.730 163.195 449.050 ;
        RECT -15.140 346.540 95.670 348.730 ;
        RECT 97.880 346.540 163.195 348.730 ;
        RECT -15.140 317.480 163.195 346.540 ;
        RECT -15.140 316.230 127.370 317.480 ;
        RECT 128.910 316.230 163.195 317.480 ;
        RECT -15.140 32.420 163.195 316.230 ;
        RECT -15.140 30.730 0.850 32.420 ;
        RECT 1.960 30.940 163.195 32.420 ;
        RECT 1.960 30.730 2.630 30.940 ;
        RECT -15.140 29.220 2.630 30.730 ;
        RECT 3.860 29.220 163.195 30.940 ;
        RECT -15.140 1.540 163.195 29.220 ;
        RECT -15.140 0.030 4.030 1.540 ;
        RECT 5.520 0.030 163.195 1.540 ;
        RECT -15.140 -1.150 163.195 0.030 ;
        RECT -15.140 -2.230 5.000 -1.150 ;
        RECT 6.490 -2.230 163.195 -1.150 ;
        RECT -15.140 -3.190 163.195 -2.230 ;
        RECT -15.140 -4.700 3.700 -3.190 ;
        RECT 5.190 -4.700 163.195 -3.190 ;
        RECT -15.140 -4.860 163.195 -4.700 ;
      LAYER met4 ;
        RECT -15.140 -4.960 163.345 482.040 ;
      LAYER met5 ;
        RECT 7.815 141.020 158.600 469.590 ;
  END
END EF_ADCS1008NC
END LIBRARY

