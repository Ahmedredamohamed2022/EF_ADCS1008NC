VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO EF_ADCS1008NC
  CLASS BLOCK ;
  FOREIGN EF_ADCS1008NC ;
  ORIGIN 16.070 4.960 ;
  SIZE 180.100 BY 489.030 ;
  PIN VSS
    ANTENNAGATEAREA 130.000000 ;
    ANTENNADIFFAREA 530.402893 ;
    PORT
      LAYER met3 ;
        RECT 96.070 346.940 97.480 348.330 ;
    END
  END VSS
  PIN HOLD
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.360000 ;
    PORT
      LAYER met3 ;
        RECT -15.970 404.980 -11.980 406.030 ;
    END
  END HOLD
  PIN EN
    ANTENNAGATEAREA 1.500000 ;
    ANTENNADIFFAREA 1.080000 ;
    PORT
      LAYER met3 ;
        RECT -16.010 383.990 -12.020 385.040 ;
    END
  END EN
  PIN DATA[9]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -15.750 316.990 -11.760 318.040 ;
    END
  END DATA[9]
  PIN DATA[8]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -15.760 281.030 -11.770 282.080 ;
    END
  END DATA[8]
  PIN DATA[7]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -16.040 250.970 -12.000 252.040 ;
    END
  END DATA[7]
  PIN DATA[6]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -16.030 218.990 -11.990 220.060 ;
    END
  END DATA[6]
  PIN DATA[5]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -16.040 183.990 -11.990 185.270 ;
    END
  END DATA[5]
  PIN DATA[4]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -16.020 151.900 -11.970 153.180 ;
    END
  END DATA[4]
  PIN DATA[3]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -16.020 117.940 -11.970 119.220 ;
    END
  END DATA[3]
  PIN DATA[2]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -16.050 83.000 -12.000 84.280 ;
    END
  END DATA[2]
  PIN DATA[1]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -16.020 48.990 -11.970 50.270 ;
    END
  END DATA[1]
  PIN VL
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met3 ;
        RECT -16.000 17.920 -11.950 19.200 ;
    END
  END VL
  PIN VH
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met3 ;
        RECT -16.030 16.030 -11.980 17.310 ;
    END
  END VH
  PIN DATA[0]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -16.020 12.850 -11.970 14.130 ;
    END
  END DATA[0]
  PIN DVDD
    ANTENNAGATEAREA 47.261497 ;
    ANTENNADIFFAREA 92.613647 ;
    PORT
      LAYER met3 ;
        RECT -16.070 0.150 -12.030 1.970 ;
    END
  END DVDD
  PIN DVSS
    ANTENNAGATEAREA 74.759102 ;
    ANTENNADIFFAREA 816.096802 ;
    PORT
      LAYER met3 ;
        RECT -16.000 -2.250 -11.960 -0.430 ;
    END
  END DVSS
  PIN VDD
    ANTENNAGATEAREA 100.000000 ;
    ANTENNADIFFAREA 2017.665894 ;
    PORT
      LAYER met3 ;
        RECT -16.020 -4.790 -11.980 -2.970 ;
    END
  END VDD
  PIN B[0]
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 160.000 449.210 163.980 450.050 ;
    END
  END B[0]
  PIN B[1]
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 160.000 447.760 163.980 448.600 ;
    END
  END B[1]
  PIN B[2]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 160.030 446.320 164.010 447.160 ;
    END
  END B[2]
  PIN CMP
    ANTENNADIFFAREA 0.492900 ;
    PORT
      LAYER met3 ;
        RECT 159.780 421.910 164.030 423.050 ;
    END
  END CMP
  PIN RST
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER met3 ;
        RECT 159.990 316.320 163.990 317.550 ;
    END
  END RST
  PIN VIN[7]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 5.760 479.990 6.730 484.010 ;
    END
  END VIN[7]
  PIN VIN[6]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 22.910 479.090 23.970 484.030 ;
    END
  END VIN[6]
  PIN VIN[5]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 39.620 479.090 40.680 484.030 ;
    END
  END VIN[5]
  PIN VIN[4]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 56.750 479.060 57.810 484.000 ;
    END
  END VIN[4]
  PIN VIN[3]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 73.500 479.090 74.560 484.030 ;
    END
  END VIN[3]
  PIN VIN[2]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 90.890 479.130 91.950 484.070 ;
    END
  END VIN[2]
  PIN VIN[1]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 107.470 479.090 108.530 484.030 ;
    END
  END VIN[1]
  PIN VIN[0]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 124.350 479.090 125.410 484.030 ;
    END
  END VIN[0]
  OBS
      LAYER li1 ;
        RECT -8.600 7.615 161.965 469.590 ;
      LAYER met1 ;
        RECT -15.720 5.090 162.120 469.590 ;
      LAYER met2 ;
        RECT -15.720 479.710 5.480 482.840 ;
        RECT 7.010 479.710 22.630 482.840 ;
        RECT -15.720 478.810 22.630 479.710 ;
        RECT 24.250 478.810 39.340 482.840 ;
        RECT 40.960 478.810 56.470 482.840 ;
        RECT -15.720 478.780 56.470 478.810 ;
        RECT 58.090 478.810 73.220 482.840 ;
        RECT 74.840 478.850 90.610 482.840 ;
        RECT 92.230 478.850 107.190 482.840 ;
        RECT 74.840 478.810 107.190 478.850 ;
        RECT 108.810 478.810 124.070 482.840 ;
        RECT 125.690 478.810 162.765 482.840 ;
        RECT 58.090 478.780 162.765 478.810 ;
        RECT -15.720 3.010 162.765 478.780 ;
      LAYER met3 ;
        RECT -16.020 450.450 163.930 482.050 ;
        RECT -16.020 447.360 159.600 450.450 ;
        RECT -16.020 445.920 159.630 447.360 ;
        RECT -16.020 423.450 163.930 445.920 ;
        RECT -16.020 421.510 159.380 423.450 ;
        RECT -16.020 406.430 163.930 421.510 ;
        RECT -11.580 404.580 163.930 406.430 ;
        RECT -16.020 385.440 163.930 404.580 ;
        RECT -11.620 383.590 163.930 385.440 ;
        RECT -16.020 348.730 163.930 383.590 ;
        RECT -16.020 346.540 95.670 348.730 ;
        RECT 97.880 346.540 163.930 348.730 ;
        RECT -16.020 318.440 163.930 346.540 ;
        RECT -11.360 317.950 163.930 318.440 ;
        RECT -11.360 316.590 159.590 317.950 ;
        RECT -16.020 315.920 159.590 316.590 ;
        RECT -16.020 282.480 163.930 315.920 ;
        RECT -11.370 280.630 163.930 282.480 ;
        RECT -16.020 252.440 163.930 280.630 ;
        RECT -11.600 250.570 163.930 252.440 ;
        RECT -16.020 220.460 163.930 250.570 ;
        RECT -11.590 218.590 163.930 220.460 ;
        RECT -16.020 185.670 163.930 218.590 ;
        RECT -11.590 183.590 163.930 185.670 ;
        RECT -16.020 153.580 163.930 183.590 ;
        RECT -11.570 151.500 163.930 153.580 ;
        RECT -16.020 119.620 163.930 151.500 ;
        RECT -11.570 117.540 163.930 119.620 ;
        RECT -16.020 84.680 163.930 117.540 ;
        RECT -11.600 82.600 163.930 84.680 ;
        RECT -16.020 50.670 163.930 82.600 ;
        RECT -11.570 48.590 163.930 50.670 ;
        RECT -16.020 19.600 163.930 48.590 ;
        RECT -11.550 17.520 163.930 19.600 ;
        RECT -11.580 15.630 163.930 17.520 ;
        RECT -16.020 14.530 163.930 15.630 ;
        RECT -11.570 12.450 163.930 14.530 ;
        RECT -16.020 2.370 163.930 12.450 ;
        RECT -11.630 -0.030 163.930 2.370 ;
        RECT -11.560 -2.650 163.930 -0.030 ;
        RECT -11.580 -4.860 163.930 -2.650 ;
      LAYER met4 ;
        RECT -15.140 -4.960 163.345 482.040 ;
      LAYER met5 ;
        RECT 7.815 141.020 158.600 469.590 ;
  END
END EF_ADCS1008NC
END LIBRARY

