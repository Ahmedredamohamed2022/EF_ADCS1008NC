magic
tech sky130A
magscale 1 2
timestamp 1694031861
<< pwell >>
rect -268 -348 268 348
<< mvnmos >>
rect -50 -100 50 100
<< mvndiff >>
rect -108 85 -50 100
rect -108 51 -96 85
rect -62 51 -50 85
rect -108 17 -50 51
rect -108 -17 -96 17
rect -62 -17 -50 17
rect -108 -51 -50 -17
rect -108 -85 -96 -51
rect -62 -85 -50 -51
rect -108 -100 -50 -85
rect 50 85 108 100
rect 50 51 62 85
rect 96 51 108 85
rect 50 17 108 51
rect 50 -17 62 17
rect 96 -17 108 17
rect 50 -51 108 -17
rect 50 -85 62 -51
rect 96 -85 108 -51
rect 50 -100 108 -85
<< mvndiffc >>
rect -96 51 -62 85
rect -96 -17 -62 17
rect -96 -85 -62 -51
rect 62 51 96 85
rect 62 -17 96 17
rect 62 -85 96 -51
<< mvpsubdiff >>
rect -242 310 242 322
rect -242 276 -119 310
rect -85 276 -51 310
rect -17 276 17 310
rect 51 276 85 310
rect 119 276 242 310
rect -242 264 242 276
rect -242 -264 -184 264
rect 184 187 242 264
rect 184 153 196 187
rect 230 153 242 187
rect 184 119 242 153
rect 184 85 196 119
rect 230 85 242 119
rect 184 51 242 85
rect 184 17 196 51
rect 230 17 242 51
rect 184 -17 242 17
rect 184 -51 196 -17
rect 230 -51 242 -17
rect 184 -85 242 -51
rect 184 -119 196 -85
rect 230 -119 242 -85
rect 184 -153 242 -119
rect 184 -187 196 -153
rect 230 -187 242 -153
rect 184 -264 242 -187
rect -242 -276 242 -264
rect -242 -310 -119 -276
rect -85 -310 -51 -276
rect -17 -310 17 -276
rect 51 -310 85 -276
rect 119 -310 242 -276
rect -242 -322 242 -310
<< mvpsubdiffcont >>
rect -119 276 -85 310
rect -51 276 -17 310
rect 17 276 51 310
rect 85 276 119 310
rect 196 153 230 187
rect 196 85 230 119
rect 196 17 230 51
rect 196 -51 230 -17
rect 196 -119 230 -85
rect 196 -187 230 -153
rect -119 -310 -85 -276
rect -51 -310 -17 -276
rect 17 -310 51 -276
rect 85 -310 119 -276
<< poly >>
rect -50 172 50 188
rect -50 138 -17 172
rect 17 138 50 172
rect -50 100 50 138
rect -50 -138 50 -100
rect -50 -172 -17 -138
rect 17 -172 50 -138
rect -50 -188 50 -172
<< polycont >>
rect -17 138 17 172
rect -17 -172 17 -138
<< locali >>
rect -230 276 -119 310
rect -85 276 -51 310
rect -17 276 17 310
rect 51 276 85 310
rect 119 276 230 310
rect -230 -276 -196 276
rect 196 187 230 276
rect -50 138 -17 172
rect 17 138 50 172
rect 196 119 230 153
rect -96 85 -62 104
rect -96 17 -62 19
rect -96 -19 -62 -17
rect -96 -104 -62 -85
rect 62 85 96 104
rect 62 17 96 19
rect 62 -19 96 -17
rect 62 -104 96 -85
rect 196 51 230 85
rect 196 -17 230 17
rect 196 -85 230 -51
rect -50 -172 -17 -138
rect 17 -172 50 -138
rect 196 -153 230 -119
rect 196 -276 230 -187
rect -230 -310 -119 -276
rect -85 -310 -51 -276
rect -17 -310 17 -276
rect 51 -310 85 -276
rect 119 -310 230 -276
<< viali >>
rect -17 138 17 172
rect -96 51 -62 53
rect -96 19 -62 51
rect -96 -51 -62 -19
rect -96 -53 -62 -51
rect 62 51 96 53
rect 62 19 96 51
rect 62 -51 96 -19
rect 62 -53 96 -51
rect -17 -172 17 -138
<< metal1 >>
rect -46 172 46 178
rect -46 138 -17 172
rect 17 138 46 172
rect -46 132 46 138
rect -102 53 -56 100
rect -102 19 -96 53
rect -62 19 -56 53
rect -102 -19 -56 19
rect -102 -53 -96 -19
rect -62 -53 -56 -19
rect -102 -100 -56 -53
rect 56 53 102 100
rect 56 19 62 53
rect 96 19 102 53
rect 56 -19 102 19
rect 56 -53 62 -19
rect 96 -53 102 -19
rect 56 -100 102 -53
rect -46 -138 46 -132
rect -46 -172 -17 -138
rect 17 -172 46 -138
rect -46 -178 46 -172
<< properties >>
string FIXED_BBOX -212 -292 212 292
<< end >>
