magic
tech sky130A
magscale 1 2
timestamp 1693827120
<< metal1 >>
rect -45300 6870 -44812 7100
rect -38676 6882 -38108 7056
rect -31876 6834 -31266 7062
rect -25268 6838 -24714 7056
rect -18430 6882 -17910 7094
rect -11268 6874 -11002 7108
rect -4764 6864 -4318 7066
rect 2000 6864 2330 7060
rect 8730 6852 9014 7052
rect 15468 6900 15800 7062
rect -18168 845 -13738 1049
rect -11262 863 -7134 1067
rect -4560 853 -696 1057
rect 2176 851 7018 1055
rect 8898 835 13148 1039
rect 15646 853 19042 1057
rect -43984 176 -43032 310
rect -37448 172 -36258 300
rect -30384 162 -29400 310
rect -23796 140 -22686 268
rect -17160 166 -16390 272
rect -9756 170 -9294 312
rect -2896 178 -2482 292
rect 3966 174 4322 290
rect 10874 166 11258 270
rect 18404 166 18736 282
<< metal3 >>
rect -18529 4687 -14255 4913
rect -8357 4715 -7847 4941
rect -1665 4713 -1146 4939
rect 5061 4697 5557 4923
rect 11805 4715 12326 4941
rect 15349 4715 19001 4941
rect -11465 1612 -4450 1622
rect -11465 1610 2162 1612
rect 8658 1610 19118 1612
rect -11465 1604 19118 1610
rect -14946 1442 19118 1604
rect -14946 1424 -11296 1442
rect -4737 1432 19118 1442
rect 1977 1430 8826 1432
rect -17685 -233 16404 -208
rect -17685 -234 15938 -233
rect -17685 -237 2453 -234
rect -17685 -257 -4229 -237
rect -17685 -401 -11000 -257
rect -10856 -381 -4229 -257
rect -4085 -378 2453 -237
rect 2597 -243 15938 -234
rect 2597 -378 9169 -243
rect -4085 -381 9169 -378
rect -10856 -387 9169 -381
rect 9313 -377 15938 -243
rect 16082 -377 16404 -233
rect 9313 -387 16404 -377
rect -10856 -401 16404 -387
rect -17685 -418 16404 -401
rect -18077 -602 15806 -600
rect -18077 -625 16400 -602
rect -18077 -633 -7579 -625
rect -18077 -777 -14332 -633
rect -14188 -769 -7579 -633
rect -7435 -633 16400 -625
rect -7435 -769 -856 -633
rect -14188 -777 -856 -769
rect -712 -635 12594 -633
rect -712 -777 5829 -635
rect -18077 -779 5829 -777
rect 5973 -777 12594 -635
rect 12738 -777 16400 -633
rect 5973 -779 16400 -777
rect -18077 -798 16400 -779
rect 12570 -800 16400 -798
<< via3 >>
rect -11000 -401 -10856 -257
rect -4229 -381 -4085 -237
rect 2453 -378 2597 -234
rect 9169 -387 9313 -243
rect 15938 -377 16082 -233
rect -14332 -777 -14188 -633
rect -7579 -769 -7435 -625
rect -856 -777 -712 -633
rect 5829 -779 5973 -635
rect 12594 -777 12738 -633
<< metal4 >>
rect -14360 -633 -14140 2974
rect -11022 -202 -10802 2966
rect -11034 -257 -10796 -202
rect -11034 -401 -11000 -257
rect -10856 -401 -10796 -257
rect -11034 -422 -10796 -401
rect -14360 -777 -14332 -633
rect -14188 -777 -14140 -633
rect -14360 -794 -14140 -777
rect -7608 -625 -7400 2970
rect -4264 -237 -4056 3372
rect -4264 -381 -4229 -237
rect -4085 -381 -4056 -237
rect -4264 -402 -4056 -381
rect -4260 -424 -4058 -402
rect -7608 -769 -7579 -625
rect -7435 -769 -7400 -625
rect -7608 -804 -7400 -769
rect -882 -633 -692 3136
rect 2422 -234 2624 3063
rect 2422 -378 2453 -234
rect 2597 -378 2624 -234
rect 2422 -415 2624 -378
rect -882 -777 -856 -633
rect -712 -777 -692 -633
rect -882 -799 -692 -777
rect 5796 -635 6008 3168
rect 9140 -243 9342 2840
rect 9140 -387 9169 -243
rect 9313 -387 9342 -243
rect 9140 -421 9342 -387
rect 5796 -779 5829 -635
rect 5973 -779 6008 -635
rect 5796 -796 6008 -779
rect 12570 -633 12766 2776
rect 15910 -233 16120 3450
rect 15910 -377 15938 -233
rect 16082 -377 16120 -233
rect 15910 -407 16120 -377
rect 12570 -777 12594 -633
rect 12738 -777 12766 -633
rect 12570 -800 12766 -777
use EF_AMUX21_ARRAY_m1  EF_AMUX21_ARRAY_m1_0
timestamp 1693827120
transform 1 0 -33884 0 1 2
box -14814 -804 19118 7108
use EF_AMUX21m  EF_AMUX21m_0
timestamp 1693827120
transform -1 0 -4821 0 1 658
box 3364 -792 9993 6424
use EF_AMUX21m  EF_AMUX21m_1
timestamp 1693827120
transform -1 0 22093 0 1 648
box 3364 -792 9993 6424
use EF_AMUX21m  EF_AMUX21m_2
timestamp 1693827120
transform -1 0 15311 0 1 630
box 3364 -792 9993 6424
use EF_AMUX21m  EF_AMUX21m_3
timestamp 1693827120
transform -1 0 8621 0 1 646
box 3364 -792 9993 6424
use EF_AMUX21m  EF_AMUX21m_4
timestamp 1693827120
transform -1 0 1907 0 1 648
box 3364 -792 9993 6424
use via14  via14_0
timestamp 1693827120
transform 1 0 -872 0 1 2788
box -14 -4 196 1202
use via14  via14_1
timestamp 1693827120
transform 1 0 15930 0 1 2734
box -14 -4 196 1202
use via14  via14_2
timestamp 1693827120
transform 1 0 12586 0 1 2760
box -14 -4 196 1202
use via14  via14_3
timestamp 1693827120
transform 1 0 9164 0 1 2732
box -14 -4 196 1202
use via14  via14_4
timestamp 1693827120
transform 1 0 5820 0 1 2756
box -14 -4 196 1202
use via14  via14_5
timestamp 1693827120
transform 1 0 2446 0 1 2768
box -14 -4 196 1202
use via14  via14_6
timestamp 1693827120
transform 1 0 -14328 0 1 2768
box -14 -4 196 1202
use via14  via14_7
timestamp 1693827120
transform 1 0 -4242 0 1 2766
box -14 -4 196 1202
use via14  via14_8
timestamp 1693827120
transform 1 0 -7594 0 1 2752
box -14 -4 196 1202
use via14  via14_9
timestamp 1693827120
transform 1 0 -10990 0 1 2740
box -14 -4 196 1202
<< labels >>
flabel metal1 s 15550 6974 15684 7034 0 FreeSans 655 0 0 0 D0
port 1 nsew
flabel metal3 s 18834 4752 18928 4910 0 FreeSans 655 0 0 0 VDD
port 2 nsew
flabel metal1 s 18852 878 18946 1006 0 FreeSans 655 0 0 0 DVSS
port 3 nsew
flabel metal1 s 18488 184 18540 242 0 FreeSans 655 0 0 0 SELD0
port 4 nsew
flabel metal3 s 14724 -380 14844 -302 0 FreeSans 655 0 0 0 VH
port 5 nsew
flabel metal3 s 13514 -746 13634 -668 0 FreeSans 655 0 0 0 VL
port 6 nsew
flabel metal1 s 11018 186 11130 248 0 FreeSans 524 0 0 0 SELD1
port 7 nsew
flabel metal1 s 8790 6892 8902 7006 0 FreeSans 524 0 0 0 D1
port 8 nsew
flabel metal3 s 18846 1472 18938 1558 0 FreeSans 524 0 0 0 DVDD
port 9 nsew
flabel metal1 s 2130 6916 2248 7002 0 FreeSans 524 0 0 0 D2
port 10 nsew
flabel metal1 s 4110 204 4224 282 0 FreeSans 524 0 0 0 SELD2
port 11 nsew
flabel metal1 s -2706 202 -2662 260 0 FreeSans 524 0 0 0 SELD3
port 12 nsew
flabel metal1 s -4570 6916 -4450 7002 0 FreeSans 524 0 0 0 D3
port 13 nsew
flabel metal1 s -9664 202 -9522 276 0 FreeSans 524 0 0 0 SELD4
port 14 nsew
flabel metal1 s -11158 6926 -11044 7012 0 FreeSans 524 0 0 0 D4
port 15 nsew
flabel metal1 s -18318 6940 -18212 6994 0 FreeSans 419 0 0 0 D5
port 16 nsew
flabel metal1 s -25066 6892 -24916 6962 0 FreeSans 419 0 0 0 D6
port 17 nsew
flabel metal1 s -31648 6876 -31520 6978 0 FreeSans 419 0 0 0 D7
port 18 nsew
flabel metal1 s -38554 6902 -38320 6998 0 FreeSans 419 0 0 0 D8
port 19 nsew
flabel metal1 s -45162 6930 -44992 7030 0 FreeSans 419 0 0 0 D9
port 20 nsew
flabel metal1 s -43776 208 -43584 284 0 FreeSans 419 0 0 0 SELD9
port 21 nsew
flabel metal1 s -30170 192 -30000 268 0 FreeSans 210 0 0 0 SELD7
port 22 nsew
flabel metal1 s -23414 162 -23322 230 0 FreeSans 210 0 0 0 SELD6
port 23 nsew
flabel metal1 s -16810 198 -16714 252 0 FreeSans 210 0 0 0 SELD5
port 24 nsew
flabel metal1 s -37126 206 -37040 272 0 FreeSans 210 0 0 0 SELD8
port 25 nsew
<< end >>
