magic
tech sky130A
magscale 1 2
timestamp 1699926577
<< metal3 >>
rect -2556 2312 2556 2340
rect -2556 2248 2472 2312
rect 2536 2248 2556 2312
rect -2556 2232 2556 2248
rect -2556 2168 2472 2232
rect 2536 2168 2556 2232
rect -2556 2152 2556 2168
rect -2556 2088 2472 2152
rect 2536 2088 2556 2152
rect -2556 2072 2556 2088
rect -2556 2008 2472 2072
rect 2536 2008 2556 2072
rect -2556 1992 2556 2008
rect -2556 1928 2472 1992
rect 2536 1928 2556 1992
rect -2556 1912 2556 1928
rect -2556 1848 2472 1912
rect 2536 1848 2556 1912
rect -2556 1832 2556 1848
rect -2556 1768 2472 1832
rect 2536 1768 2556 1832
rect -2556 1752 2556 1768
rect -2556 1688 2472 1752
rect 2536 1688 2556 1752
rect -2556 1672 2556 1688
rect -2556 1608 2472 1672
rect 2536 1608 2556 1672
rect -2556 1592 2556 1608
rect -2556 1528 2472 1592
rect 2536 1528 2556 1592
rect -2556 1512 2556 1528
rect -2556 1448 2472 1512
rect 2536 1448 2556 1512
rect -2556 1432 2556 1448
rect -2556 1368 2472 1432
rect 2536 1368 2556 1432
rect -2556 1352 2556 1368
rect -2556 1288 2472 1352
rect 2536 1288 2556 1352
rect -2556 1272 2556 1288
rect -2556 1208 2472 1272
rect 2536 1208 2556 1272
rect -2556 1192 2556 1208
rect -2556 1128 2472 1192
rect 2536 1128 2556 1192
rect -2556 1112 2556 1128
rect -2556 1048 2472 1112
rect 2536 1048 2556 1112
rect -2556 1032 2556 1048
rect -2556 968 2472 1032
rect 2536 968 2556 1032
rect -2556 952 2556 968
rect -2556 888 2472 952
rect 2536 888 2556 952
rect -2556 872 2556 888
rect -2556 808 2472 872
rect 2536 808 2556 872
rect -2556 792 2556 808
rect -2556 728 2472 792
rect 2536 728 2556 792
rect -2556 712 2556 728
rect -2556 648 2472 712
rect 2536 648 2556 712
rect -2556 632 2556 648
rect -2556 568 2472 632
rect 2536 568 2556 632
rect -2556 552 2556 568
rect -2556 488 2472 552
rect 2536 488 2556 552
rect -2556 472 2556 488
rect -2556 408 2472 472
rect 2536 408 2556 472
rect -2556 392 2556 408
rect -2556 328 2472 392
rect 2536 328 2556 392
rect -2556 312 2556 328
rect -2556 248 2472 312
rect 2536 248 2556 312
rect -2556 232 2556 248
rect -2556 168 2472 232
rect 2536 168 2556 232
rect -2556 152 2556 168
rect -2556 88 2472 152
rect 2536 88 2556 152
rect -2556 72 2556 88
rect -2556 8 2472 72
rect 2536 8 2556 72
rect -2556 -8 2556 8
rect -2556 -72 2472 -8
rect 2536 -72 2556 -8
rect -2556 -88 2556 -72
rect -2556 -152 2472 -88
rect 2536 -152 2556 -88
rect -2556 -168 2556 -152
rect -2556 -232 2472 -168
rect 2536 -232 2556 -168
rect -2556 -248 2556 -232
rect -2556 -312 2472 -248
rect 2536 -312 2556 -248
rect -2556 -328 2556 -312
rect -2556 -392 2472 -328
rect 2536 -392 2556 -328
rect -2556 -408 2556 -392
rect -2556 -472 2472 -408
rect 2536 -472 2556 -408
rect -2556 -488 2556 -472
rect -2556 -552 2472 -488
rect 2536 -552 2556 -488
rect -2556 -568 2556 -552
rect -2556 -632 2472 -568
rect 2536 -632 2556 -568
rect -2556 -648 2556 -632
rect -2556 -712 2472 -648
rect 2536 -712 2556 -648
rect -2556 -728 2556 -712
rect -2556 -792 2472 -728
rect 2536 -792 2556 -728
rect -2556 -808 2556 -792
rect -2556 -872 2472 -808
rect 2536 -872 2556 -808
rect -2556 -888 2556 -872
rect -2556 -952 2472 -888
rect 2536 -952 2556 -888
rect -2556 -968 2556 -952
rect -2556 -1032 2472 -968
rect 2536 -1032 2556 -968
rect -2556 -1048 2556 -1032
rect -2556 -1112 2472 -1048
rect 2536 -1112 2556 -1048
rect -2556 -1128 2556 -1112
rect -2556 -1192 2472 -1128
rect 2536 -1192 2556 -1128
rect -2556 -1208 2556 -1192
rect -2556 -1272 2472 -1208
rect 2536 -1272 2556 -1208
rect -2556 -1288 2556 -1272
rect -2556 -1352 2472 -1288
rect 2536 -1352 2556 -1288
rect -2556 -1368 2556 -1352
rect -2556 -1432 2472 -1368
rect 2536 -1432 2556 -1368
rect -2556 -1448 2556 -1432
rect -2556 -1512 2472 -1448
rect 2536 -1512 2556 -1448
rect -2556 -1528 2556 -1512
rect -2556 -1592 2472 -1528
rect 2536 -1592 2556 -1528
rect -2556 -1608 2556 -1592
rect -2556 -1672 2472 -1608
rect 2536 -1672 2556 -1608
rect -2556 -1688 2556 -1672
rect -2556 -1752 2472 -1688
rect 2536 -1752 2556 -1688
rect -2556 -1768 2556 -1752
rect -2556 -1832 2472 -1768
rect 2536 -1832 2556 -1768
rect -2556 -1848 2556 -1832
rect -2556 -1912 2472 -1848
rect 2536 -1912 2556 -1848
rect -2556 -1928 2556 -1912
rect -2556 -1992 2472 -1928
rect 2536 -1992 2556 -1928
rect -2556 -2008 2556 -1992
rect -2556 -2072 2472 -2008
rect 2536 -2072 2556 -2008
rect -2556 -2088 2556 -2072
rect -2556 -2152 2472 -2088
rect 2536 -2152 2556 -2088
rect -2556 -2168 2556 -2152
rect -2556 -2232 2472 -2168
rect 2536 -2232 2556 -2168
rect -2556 -2248 2556 -2232
rect -2556 -2312 2472 -2248
rect 2536 -2312 2556 -2248
rect -2556 -2340 2556 -2312
<< via3 >>
rect 2472 2248 2536 2312
rect 2472 2168 2536 2232
rect 2472 2088 2536 2152
rect 2472 2008 2536 2072
rect 2472 1928 2536 1992
rect 2472 1848 2536 1912
rect 2472 1768 2536 1832
rect 2472 1688 2536 1752
rect 2472 1608 2536 1672
rect 2472 1528 2536 1592
rect 2472 1448 2536 1512
rect 2472 1368 2536 1432
rect 2472 1288 2536 1352
rect 2472 1208 2536 1272
rect 2472 1128 2536 1192
rect 2472 1048 2536 1112
rect 2472 968 2536 1032
rect 2472 888 2536 952
rect 2472 808 2536 872
rect 2472 728 2536 792
rect 2472 648 2536 712
rect 2472 568 2536 632
rect 2472 488 2536 552
rect 2472 408 2536 472
rect 2472 328 2536 392
rect 2472 248 2536 312
rect 2472 168 2536 232
rect 2472 88 2536 152
rect 2472 8 2536 72
rect 2472 -72 2536 -8
rect 2472 -152 2536 -88
rect 2472 -232 2536 -168
rect 2472 -312 2536 -248
rect 2472 -392 2536 -328
rect 2472 -472 2536 -408
rect 2472 -552 2536 -488
rect 2472 -632 2536 -568
rect 2472 -712 2536 -648
rect 2472 -792 2536 -728
rect 2472 -872 2536 -808
rect 2472 -952 2536 -888
rect 2472 -1032 2536 -968
rect 2472 -1112 2536 -1048
rect 2472 -1192 2536 -1128
rect 2472 -1272 2536 -1208
rect 2472 -1352 2536 -1288
rect 2472 -1432 2536 -1368
rect 2472 -1512 2536 -1448
rect 2472 -1592 2536 -1528
rect 2472 -1672 2536 -1608
rect 2472 -1752 2536 -1688
rect 2472 -1832 2536 -1768
rect 2472 -1912 2536 -1848
rect 2472 -1992 2536 -1928
rect 2472 -2072 2536 -2008
rect 2472 -2152 2536 -2088
rect 2472 -2232 2536 -2168
rect 2472 -2312 2536 -2248
<< mimcap >>
rect -2516 2232 2224 2300
rect -2516 -2232 -2458 2232
rect 2166 -2232 2224 2232
rect -2516 -2300 2224 -2232
<< mimcapcontact >>
rect -2458 -2232 2166 2232
<< metal4 >>
rect 2456 2312 2552 2328
rect -2477 2232 2185 2261
rect -2477 -2232 -2458 2232
rect 2166 -2232 2185 2232
rect -2477 -2261 2185 -2232
rect 2456 2248 2472 2312
rect 2536 2248 2552 2312
rect 2456 2232 2552 2248
rect 2456 2168 2472 2232
rect 2536 2168 2552 2232
rect 2456 2152 2552 2168
rect 2456 2088 2472 2152
rect 2536 2088 2552 2152
rect 2456 2072 2552 2088
rect 2456 2008 2472 2072
rect 2536 2008 2552 2072
rect 2456 1992 2552 2008
rect 2456 1928 2472 1992
rect 2536 1928 2552 1992
rect 2456 1912 2552 1928
rect 2456 1848 2472 1912
rect 2536 1848 2552 1912
rect 2456 1832 2552 1848
rect 2456 1768 2472 1832
rect 2536 1768 2552 1832
rect 2456 1752 2552 1768
rect 2456 1688 2472 1752
rect 2536 1688 2552 1752
rect 2456 1672 2552 1688
rect 2456 1608 2472 1672
rect 2536 1608 2552 1672
rect 2456 1592 2552 1608
rect 2456 1528 2472 1592
rect 2536 1528 2552 1592
rect 2456 1512 2552 1528
rect 2456 1448 2472 1512
rect 2536 1448 2552 1512
rect 2456 1432 2552 1448
rect 2456 1368 2472 1432
rect 2536 1368 2552 1432
rect 2456 1352 2552 1368
rect 2456 1288 2472 1352
rect 2536 1288 2552 1352
rect 2456 1272 2552 1288
rect 2456 1208 2472 1272
rect 2536 1208 2552 1272
rect 2456 1192 2552 1208
rect 2456 1128 2472 1192
rect 2536 1128 2552 1192
rect 2456 1112 2552 1128
rect 2456 1048 2472 1112
rect 2536 1048 2552 1112
rect 2456 1032 2552 1048
rect 2456 968 2472 1032
rect 2536 968 2552 1032
rect 2456 952 2552 968
rect 2456 888 2472 952
rect 2536 888 2552 952
rect 2456 872 2552 888
rect 2456 808 2472 872
rect 2536 808 2552 872
rect 2456 792 2552 808
rect 2456 728 2472 792
rect 2536 728 2552 792
rect 2456 712 2552 728
rect 2456 648 2472 712
rect 2536 648 2552 712
rect 2456 632 2552 648
rect 2456 568 2472 632
rect 2536 568 2552 632
rect 2456 552 2552 568
rect 2456 488 2472 552
rect 2536 488 2552 552
rect 2456 472 2552 488
rect 2456 408 2472 472
rect 2536 408 2552 472
rect 2456 392 2552 408
rect 2456 328 2472 392
rect 2536 328 2552 392
rect 2456 312 2552 328
rect 2456 248 2472 312
rect 2536 248 2552 312
rect 2456 232 2552 248
rect 2456 168 2472 232
rect 2536 168 2552 232
rect 2456 152 2552 168
rect 2456 88 2472 152
rect 2536 88 2552 152
rect 2456 72 2552 88
rect 2456 8 2472 72
rect 2536 8 2552 72
rect 2456 -8 2552 8
rect 2456 -72 2472 -8
rect 2536 -72 2552 -8
rect 2456 -88 2552 -72
rect 2456 -152 2472 -88
rect 2536 -152 2552 -88
rect 2456 -168 2552 -152
rect 2456 -232 2472 -168
rect 2536 -232 2552 -168
rect 2456 -248 2552 -232
rect 2456 -312 2472 -248
rect 2536 -312 2552 -248
rect 2456 -328 2552 -312
rect 2456 -392 2472 -328
rect 2536 -392 2552 -328
rect 2456 -408 2552 -392
rect 2456 -472 2472 -408
rect 2536 -472 2552 -408
rect 2456 -488 2552 -472
rect 2456 -552 2472 -488
rect 2536 -552 2552 -488
rect 2456 -568 2552 -552
rect 2456 -632 2472 -568
rect 2536 -632 2552 -568
rect 2456 -648 2552 -632
rect 2456 -712 2472 -648
rect 2536 -712 2552 -648
rect 2456 -728 2552 -712
rect 2456 -792 2472 -728
rect 2536 -792 2552 -728
rect 2456 -808 2552 -792
rect 2456 -872 2472 -808
rect 2536 -872 2552 -808
rect 2456 -888 2552 -872
rect 2456 -952 2472 -888
rect 2536 -952 2552 -888
rect 2456 -968 2552 -952
rect 2456 -1032 2472 -968
rect 2536 -1032 2552 -968
rect 2456 -1048 2552 -1032
rect 2456 -1112 2472 -1048
rect 2536 -1112 2552 -1048
rect 2456 -1128 2552 -1112
rect 2456 -1192 2472 -1128
rect 2536 -1192 2552 -1128
rect 2456 -1208 2552 -1192
rect 2456 -1272 2472 -1208
rect 2536 -1272 2552 -1208
rect 2456 -1288 2552 -1272
rect 2456 -1352 2472 -1288
rect 2536 -1352 2552 -1288
rect 2456 -1368 2552 -1352
rect 2456 -1432 2472 -1368
rect 2536 -1432 2552 -1368
rect 2456 -1448 2552 -1432
rect 2456 -1512 2472 -1448
rect 2536 -1512 2552 -1448
rect 2456 -1528 2552 -1512
rect 2456 -1592 2472 -1528
rect 2536 -1592 2552 -1528
rect 2456 -1608 2552 -1592
rect 2456 -1672 2472 -1608
rect 2536 -1672 2552 -1608
rect 2456 -1688 2552 -1672
rect 2456 -1752 2472 -1688
rect 2536 -1752 2552 -1688
rect 2456 -1768 2552 -1752
rect 2456 -1832 2472 -1768
rect 2536 -1832 2552 -1768
rect 2456 -1848 2552 -1832
rect 2456 -1912 2472 -1848
rect 2536 -1912 2552 -1848
rect 2456 -1928 2552 -1912
rect 2456 -1992 2472 -1928
rect 2536 -1992 2552 -1928
rect 2456 -2008 2552 -1992
rect 2456 -2072 2472 -2008
rect 2536 -2072 2552 -2008
rect 2456 -2088 2552 -2072
rect 2456 -2152 2472 -2088
rect 2536 -2152 2552 -2088
rect 2456 -2168 2552 -2152
rect 2456 -2232 2472 -2168
rect 2536 -2232 2552 -2168
rect 2456 -2248 2552 -2232
rect 2456 -2312 2472 -2248
rect 2536 -2312 2552 -2248
rect 2456 -2328 2552 -2312
<< properties >>
string FIXED_BBOX -2556 -2340 2264 2340
<< end >>
