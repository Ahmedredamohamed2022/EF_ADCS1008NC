magic
tech sky130A
magscale 1 2
timestamp 1693827120
<< nwell >>
rect -3389 -1269 3389 1269
<< mvpmos >>
rect -3131 772 -3031 972
rect -2973 772 -2873 972
rect -2815 772 -2715 972
rect -2657 772 -2557 972
rect -2499 772 -2399 972
rect -2341 772 -2241 972
rect -2183 772 -2083 972
rect -2025 772 -1925 972
rect -1867 772 -1767 972
rect -1709 772 -1609 972
rect -1551 772 -1451 972
rect -1393 772 -1293 972
rect -1235 772 -1135 972
rect -1077 772 -977 972
rect -919 772 -819 972
rect -761 772 -661 972
rect -603 772 -503 972
rect -445 772 -345 972
rect -287 772 -187 972
rect -129 772 -29 972
rect 29 772 129 972
rect 187 772 287 972
rect 345 772 445 972
rect 503 772 603 972
rect 661 772 761 972
rect 819 772 919 972
rect 977 772 1077 972
rect 1135 772 1235 972
rect 1293 772 1393 972
rect 1451 772 1551 972
rect 1609 772 1709 972
rect 1767 772 1867 972
rect 1925 772 2025 972
rect 2083 772 2183 972
rect 2241 772 2341 972
rect 2399 772 2499 972
rect 2557 772 2657 972
rect 2715 772 2815 972
rect 2873 772 2973 972
rect 3031 772 3131 972
rect -3131 336 -3031 536
rect -2973 336 -2873 536
rect -2815 336 -2715 536
rect -2657 336 -2557 536
rect -2499 336 -2399 536
rect -2341 336 -2241 536
rect -2183 336 -2083 536
rect -2025 336 -1925 536
rect -1867 336 -1767 536
rect -1709 336 -1609 536
rect -1551 336 -1451 536
rect -1393 336 -1293 536
rect -1235 336 -1135 536
rect -1077 336 -977 536
rect -919 336 -819 536
rect -761 336 -661 536
rect -603 336 -503 536
rect -445 336 -345 536
rect -287 336 -187 536
rect -129 336 -29 536
rect 29 336 129 536
rect 187 336 287 536
rect 345 336 445 536
rect 503 336 603 536
rect 661 336 761 536
rect 819 336 919 536
rect 977 336 1077 536
rect 1135 336 1235 536
rect 1293 336 1393 536
rect 1451 336 1551 536
rect 1609 336 1709 536
rect 1767 336 1867 536
rect 1925 336 2025 536
rect 2083 336 2183 536
rect 2241 336 2341 536
rect 2399 336 2499 536
rect 2557 336 2657 536
rect 2715 336 2815 536
rect 2873 336 2973 536
rect 3031 336 3131 536
rect -3131 -100 -3031 100
rect -2973 -100 -2873 100
rect -2815 -100 -2715 100
rect -2657 -100 -2557 100
rect -2499 -100 -2399 100
rect -2341 -100 -2241 100
rect -2183 -100 -2083 100
rect -2025 -100 -1925 100
rect -1867 -100 -1767 100
rect -1709 -100 -1609 100
rect -1551 -100 -1451 100
rect -1393 -100 -1293 100
rect -1235 -100 -1135 100
rect -1077 -100 -977 100
rect -919 -100 -819 100
rect -761 -100 -661 100
rect -603 -100 -503 100
rect -445 -100 -345 100
rect -287 -100 -187 100
rect -129 -100 -29 100
rect 29 -100 129 100
rect 187 -100 287 100
rect 345 -100 445 100
rect 503 -100 603 100
rect 661 -100 761 100
rect 819 -100 919 100
rect 977 -100 1077 100
rect 1135 -100 1235 100
rect 1293 -100 1393 100
rect 1451 -100 1551 100
rect 1609 -100 1709 100
rect 1767 -100 1867 100
rect 1925 -100 2025 100
rect 2083 -100 2183 100
rect 2241 -100 2341 100
rect 2399 -100 2499 100
rect 2557 -100 2657 100
rect 2715 -100 2815 100
rect 2873 -100 2973 100
rect 3031 -100 3131 100
rect -3131 -536 -3031 -336
rect -2973 -536 -2873 -336
rect -2815 -536 -2715 -336
rect -2657 -536 -2557 -336
rect -2499 -536 -2399 -336
rect -2341 -536 -2241 -336
rect -2183 -536 -2083 -336
rect -2025 -536 -1925 -336
rect -1867 -536 -1767 -336
rect -1709 -536 -1609 -336
rect -1551 -536 -1451 -336
rect -1393 -536 -1293 -336
rect -1235 -536 -1135 -336
rect -1077 -536 -977 -336
rect -919 -536 -819 -336
rect -761 -536 -661 -336
rect -603 -536 -503 -336
rect -445 -536 -345 -336
rect -287 -536 -187 -336
rect -129 -536 -29 -336
rect 29 -536 129 -336
rect 187 -536 287 -336
rect 345 -536 445 -336
rect 503 -536 603 -336
rect 661 -536 761 -336
rect 819 -536 919 -336
rect 977 -536 1077 -336
rect 1135 -536 1235 -336
rect 1293 -536 1393 -336
rect 1451 -536 1551 -336
rect 1609 -536 1709 -336
rect 1767 -536 1867 -336
rect 1925 -536 2025 -336
rect 2083 -536 2183 -336
rect 2241 -536 2341 -336
rect 2399 -536 2499 -336
rect 2557 -536 2657 -336
rect 2715 -536 2815 -336
rect 2873 -536 2973 -336
rect 3031 -536 3131 -336
rect -3131 -972 -3031 -772
rect -2973 -972 -2873 -772
rect -2815 -972 -2715 -772
rect -2657 -972 -2557 -772
rect -2499 -972 -2399 -772
rect -2341 -972 -2241 -772
rect -2183 -972 -2083 -772
rect -2025 -972 -1925 -772
rect -1867 -972 -1767 -772
rect -1709 -972 -1609 -772
rect -1551 -972 -1451 -772
rect -1393 -972 -1293 -772
rect -1235 -972 -1135 -772
rect -1077 -972 -977 -772
rect -919 -972 -819 -772
rect -761 -972 -661 -772
rect -603 -972 -503 -772
rect -445 -972 -345 -772
rect -287 -972 -187 -772
rect -129 -972 -29 -772
rect 29 -972 129 -772
rect 187 -972 287 -772
rect 345 -972 445 -772
rect 503 -972 603 -772
rect 661 -972 761 -772
rect 819 -972 919 -772
rect 977 -972 1077 -772
rect 1135 -972 1235 -772
rect 1293 -972 1393 -772
rect 1451 -972 1551 -772
rect 1609 -972 1709 -772
rect 1767 -972 1867 -772
rect 1925 -972 2025 -772
rect 2083 -972 2183 -772
rect 2241 -972 2341 -772
rect 2399 -972 2499 -772
rect 2557 -972 2657 -772
rect 2715 -972 2815 -772
rect 2873 -972 2973 -772
rect 3031 -972 3131 -772
<< mvpdiff >>
rect -3189 957 -3131 972
rect -3189 923 -3177 957
rect -3143 923 -3131 957
rect -3189 889 -3131 923
rect -3189 855 -3177 889
rect -3143 855 -3131 889
rect -3189 821 -3131 855
rect -3189 787 -3177 821
rect -3143 787 -3131 821
rect -3189 772 -3131 787
rect -3031 957 -2973 972
rect -3031 923 -3019 957
rect -2985 923 -2973 957
rect -3031 889 -2973 923
rect -3031 855 -3019 889
rect -2985 855 -2973 889
rect -3031 821 -2973 855
rect -3031 787 -3019 821
rect -2985 787 -2973 821
rect -3031 772 -2973 787
rect -2873 957 -2815 972
rect -2873 923 -2861 957
rect -2827 923 -2815 957
rect -2873 889 -2815 923
rect -2873 855 -2861 889
rect -2827 855 -2815 889
rect -2873 821 -2815 855
rect -2873 787 -2861 821
rect -2827 787 -2815 821
rect -2873 772 -2815 787
rect -2715 957 -2657 972
rect -2715 923 -2703 957
rect -2669 923 -2657 957
rect -2715 889 -2657 923
rect -2715 855 -2703 889
rect -2669 855 -2657 889
rect -2715 821 -2657 855
rect -2715 787 -2703 821
rect -2669 787 -2657 821
rect -2715 772 -2657 787
rect -2557 957 -2499 972
rect -2557 923 -2545 957
rect -2511 923 -2499 957
rect -2557 889 -2499 923
rect -2557 855 -2545 889
rect -2511 855 -2499 889
rect -2557 821 -2499 855
rect -2557 787 -2545 821
rect -2511 787 -2499 821
rect -2557 772 -2499 787
rect -2399 957 -2341 972
rect -2399 923 -2387 957
rect -2353 923 -2341 957
rect -2399 889 -2341 923
rect -2399 855 -2387 889
rect -2353 855 -2341 889
rect -2399 821 -2341 855
rect -2399 787 -2387 821
rect -2353 787 -2341 821
rect -2399 772 -2341 787
rect -2241 957 -2183 972
rect -2241 923 -2229 957
rect -2195 923 -2183 957
rect -2241 889 -2183 923
rect -2241 855 -2229 889
rect -2195 855 -2183 889
rect -2241 821 -2183 855
rect -2241 787 -2229 821
rect -2195 787 -2183 821
rect -2241 772 -2183 787
rect -2083 957 -2025 972
rect -2083 923 -2071 957
rect -2037 923 -2025 957
rect -2083 889 -2025 923
rect -2083 855 -2071 889
rect -2037 855 -2025 889
rect -2083 821 -2025 855
rect -2083 787 -2071 821
rect -2037 787 -2025 821
rect -2083 772 -2025 787
rect -1925 957 -1867 972
rect -1925 923 -1913 957
rect -1879 923 -1867 957
rect -1925 889 -1867 923
rect -1925 855 -1913 889
rect -1879 855 -1867 889
rect -1925 821 -1867 855
rect -1925 787 -1913 821
rect -1879 787 -1867 821
rect -1925 772 -1867 787
rect -1767 957 -1709 972
rect -1767 923 -1755 957
rect -1721 923 -1709 957
rect -1767 889 -1709 923
rect -1767 855 -1755 889
rect -1721 855 -1709 889
rect -1767 821 -1709 855
rect -1767 787 -1755 821
rect -1721 787 -1709 821
rect -1767 772 -1709 787
rect -1609 957 -1551 972
rect -1609 923 -1597 957
rect -1563 923 -1551 957
rect -1609 889 -1551 923
rect -1609 855 -1597 889
rect -1563 855 -1551 889
rect -1609 821 -1551 855
rect -1609 787 -1597 821
rect -1563 787 -1551 821
rect -1609 772 -1551 787
rect -1451 957 -1393 972
rect -1451 923 -1439 957
rect -1405 923 -1393 957
rect -1451 889 -1393 923
rect -1451 855 -1439 889
rect -1405 855 -1393 889
rect -1451 821 -1393 855
rect -1451 787 -1439 821
rect -1405 787 -1393 821
rect -1451 772 -1393 787
rect -1293 957 -1235 972
rect -1293 923 -1281 957
rect -1247 923 -1235 957
rect -1293 889 -1235 923
rect -1293 855 -1281 889
rect -1247 855 -1235 889
rect -1293 821 -1235 855
rect -1293 787 -1281 821
rect -1247 787 -1235 821
rect -1293 772 -1235 787
rect -1135 957 -1077 972
rect -1135 923 -1123 957
rect -1089 923 -1077 957
rect -1135 889 -1077 923
rect -1135 855 -1123 889
rect -1089 855 -1077 889
rect -1135 821 -1077 855
rect -1135 787 -1123 821
rect -1089 787 -1077 821
rect -1135 772 -1077 787
rect -977 957 -919 972
rect -977 923 -965 957
rect -931 923 -919 957
rect -977 889 -919 923
rect -977 855 -965 889
rect -931 855 -919 889
rect -977 821 -919 855
rect -977 787 -965 821
rect -931 787 -919 821
rect -977 772 -919 787
rect -819 957 -761 972
rect -819 923 -807 957
rect -773 923 -761 957
rect -819 889 -761 923
rect -819 855 -807 889
rect -773 855 -761 889
rect -819 821 -761 855
rect -819 787 -807 821
rect -773 787 -761 821
rect -819 772 -761 787
rect -661 957 -603 972
rect -661 923 -649 957
rect -615 923 -603 957
rect -661 889 -603 923
rect -661 855 -649 889
rect -615 855 -603 889
rect -661 821 -603 855
rect -661 787 -649 821
rect -615 787 -603 821
rect -661 772 -603 787
rect -503 957 -445 972
rect -503 923 -491 957
rect -457 923 -445 957
rect -503 889 -445 923
rect -503 855 -491 889
rect -457 855 -445 889
rect -503 821 -445 855
rect -503 787 -491 821
rect -457 787 -445 821
rect -503 772 -445 787
rect -345 957 -287 972
rect -345 923 -333 957
rect -299 923 -287 957
rect -345 889 -287 923
rect -345 855 -333 889
rect -299 855 -287 889
rect -345 821 -287 855
rect -345 787 -333 821
rect -299 787 -287 821
rect -345 772 -287 787
rect -187 957 -129 972
rect -187 923 -175 957
rect -141 923 -129 957
rect -187 889 -129 923
rect -187 855 -175 889
rect -141 855 -129 889
rect -187 821 -129 855
rect -187 787 -175 821
rect -141 787 -129 821
rect -187 772 -129 787
rect -29 957 29 972
rect -29 923 -17 957
rect 17 923 29 957
rect -29 889 29 923
rect -29 855 -17 889
rect 17 855 29 889
rect -29 821 29 855
rect -29 787 -17 821
rect 17 787 29 821
rect -29 772 29 787
rect 129 957 187 972
rect 129 923 141 957
rect 175 923 187 957
rect 129 889 187 923
rect 129 855 141 889
rect 175 855 187 889
rect 129 821 187 855
rect 129 787 141 821
rect 175 787 187 821
rect 129 772 187 787
rect 287 957 345 972
rect 287 923 299 957
rect 333 923 345 957
rect 287 889 345 923
rect 287 855 299 889
rect 333 855 345 889
rect 287 821 345 855
rect 287 787 299 821
rect 333 787 345 821
rect 287 772 345 787
rect 445 957 503 972
rect 445 923 457 957
rect 491 923 503 957
rect 445 889 503 923
rect 445 855 457 889
rect 491 855 503 889
rect 445 821 503 855
rect 445 787 457 821
rect 491 787 503 821
rect 445 772 503 787
rect 603 957 661 972
rect 603 923 615 957
rect 649 923 661 957
rect 603 889 661 923
rect 603 855 615 889
rect 649 855 661 889
rect 603 821 661 855
rect 603 787 615 821
rect 649 787 661 821
rect 603 772 661 787
rect 761 957 819 972
rect 761 923 773 957
rect 807 923 819 957
rect 761 889 819 923
rect 761 855 773 889
rect 807 855 819 889
rect 761 821 819 855
rect 761 787 773 821
rect 807 787 819 821
rect 761 772 819 787
rect 919 957 977 972
rect 919 923 931 957
rect 965 923 977 957
rect 919 889 977 923
rect 919 855 931 889
rect 965 855 977 889
rect 919 821 977 855
rect 919 787 931 821
rect 965 787 977 821
rect 919 772 977 787
rect 1077 957 1135 972
rect 1077 923 1089 957
rect 1123 923 1135 957
rect 1077 889 1135 923
rect 1077 855 1089 889
rect 1123 855 1135 889
rect 1077 821 1135 855
rect 1077 787 1089 821
rect 1123 787 1135 821
rect 1077 772 1135 787
rect 1235 957 1293 972
rect 1235 923 1247 957
rect 1281 923 1293 957
rect 1235 889 1293 923
rect 1235 855 1247 889
rect 1281 855 1293 889
rect 1235 821 1293 855
rect 1235 787 1247 821
rect 1281 787 1293 821
rect 1235 772 1293 787
rect 1393 957 1451 972
rect 1393 923 1405 957
rect 1439 923 1451 957
rect 1393 889 1451 923
rect 1393 855 1405 889
rect 1439 855 1451 889
rect 1393 821 1451 855
rect 1393 787 1405 821
rect 1439 787 1451 821
rect 1393 772 1451 787
rect 1551 957 1609 972
rect 1551 923 1563 957
rect 1597 923 1609 957
rect 1551 889 1609 923
rect 1551 855 1563 889
rect 1597 855 1609 889
rect 1551 821 1609 855
rect 1551 787 1563 821
rect 1597 787 1609 821
rect 1551 772 1609 787
rect 1709 957 1767 972
rect 1709 923 1721 957
rect 1755 923 1767 957
rect 1709 889 1767 923
rect 1709 855 1721 889
rect 1755 855 1767 889
rect 1709 821 1767 855
rect 1709 787 1721 821
rect 1755 787 1767 821
rect 1709 772 1767 787
rect 1867 957 1925 972
rect 1867 923 1879 957
rect 1913 923 1925 957
rect 1867 889 1925 923
rect 1867 855 1879 889
rect 1913 855 1925 889
rect 1867 821 1925 855
rect 1867 787 1879 821
rect 1913 787 1925 821
rect 1867 772 1925 787
rect 2025 957 2083 972
rect 2025 923 2037 957
rect 2071 923 2083 957
rect 2025 889 2083 923
rect 2025 855 2037 889
rect 2071 855 2083 889
rect 2025 821 2083 855
rect 2025 787 2037 821
rect 2071 787 2083 821
rect 2025 772 2083 787
rect 2183 957 2241 972
rect 2183 923 2195 957
rect 2229 923 2241 957
rect 2183 889 2241 923
rect 2183 855 2195 889
rect 2229 855 2241 889
rect 2183 821 2241 855
rect 2183 787 2195 821
rect 2229 787 2241 821
rect 2183 772 2241 787
rect 2341 957 2399 972
rect 2341 923 2353 957
rect 2387 923 2399 957
rect 2341 889 2399 923
rect 2341 855 2353 889
rect 2387 855 2399 889
rect 2341 821 2399 855
rect 2341 787 2353 821
rect 2387 787 2399 821
rect 2341 772 2399 787
rect 2499 957 2557 972
rect 2499 923 2511 957
rect 2545 923 2557 957
rect 2499 889 2557 923
rect 2499 855 2511 889
rect 2545 855 2557 889
rect 2499 821 2557 855
rect 2499 787 2511 821
rect 2545 787 2557 821
rect 2499 772 2557 787
rect 2657 957 2715 972
rect 2657 923 2669 957
rect 2703 923 2715 957
rect 2657 889 2715 923
rect 2657 855 2669 889
rect 2703 855 2715 889
rect 2657 821 2715 855
rect 2657 787 2669 821
rect 2703 787 2715 821
rect 2657 772 2715 787
rect 2815 957 2873 972
rect 2815 923 2827 957
rect 2861 923 2873 957
rect 2815 889 2873 923
rect 2815 855 2827 889
rect 2861 855 2873 889
rect 2815 821 2873 855
rect 2815 787 2827 821
rect 2861 787 2873 821
rect 2815 772 2873 787
rect 2973 957 3031 972
rect 2973 923 2985 957
rect 3019 923 3031 957
rect 2973 889 3031 923
rect 2973 855 2985 889
rect 3019 855 3031 889
rect 2973 821 3031 855
rect 2973 787 2985 821
rect 3019 787 3031 821
rect 2973 772 3031 787
rect 3131 957 3189 972
rect 3131 923 3143 957
rect 3177 923 3189 957
rect 3131 889 3189 923
rect 3131 855 3143 889
rect 3177 855 3189 889
rect 3131 821 3189 855
rect 3131 787 3143 821
rect 3177 787 3189 821
rect 3131 772 3189 787
rect -3189 521 -3131 536
rect -3189 487 -3177 521
rect -3143 487 -3131 521
rect -3189 453 -3131 487
rect -3189 419 -3177 453
rect -3143 419 -3131 453
rect -3189 385 -3131 419
rect -3189 351 -3177 385
rect -3143 351 -3131 385
rect -3189 336 -3131 351
rect -3031 521 -2973 536
rect -3031 487 -3019 521
rect -2985 487 -2973 521
rect -3031 453 -2973 487
rect -3031 419 -3019 453
rect -2985 419 -2973 453
rect -3031 385 -2973 419
rect -3031 351 -3019 385
rect -2985 351 -2973 385
rect -3031 336 -2973 351
rect -2873 521 -2815 536
rect -2873 487 -2861 521
rect -2827 487 -2815 521
rect -2873 453 -2815 487
rect -2873 419 -2861 453
rect -2827 419 -2815 453
rect -2873 385 -2815 419
rect -2873 351 -2861 385
rect -2827 351 -2815 385
rect -2873 336 -2815 351
rect -2715 521 -2657 536
rect -2715 487 -2703 521
rect -2669 487 -2657 521
rect -2715 453 -2657 487
rect -2715 419 -2703 453
rect -2669 419 -2657 453
rect -2715 385 -2657 419
rect -2715 351 -2703 385
rect -2669 351 -2657 385
rect -2715 336 -2657 351
rect -2557 521 -2499 536
rect -2557 487 -2545 521
rect -2511 487 -2499 521
rect -2557 453 -2499 487
rect -2557 419 -2545 453
rect -2511 419 -2499 453
rect -2557 385 -2499 419
rect -2557 351 -2545 385
rect -2511 351 -2499 385
rect -2557 336 -2499 351
rect -2399 521 -2341 536
rect -2399 487 -2387 521
rect -2353 487 -2341 521
rect -2399 453 -2341 487
rect -2399 419 -2387 453
rect -2353 419 -2341 453
rect -2399 385 -2341 419
rect -2399 351 -2387 385
rect -2353 351 -2341 385
rect -2399 336 -2341 351
rect -2241 521 -2183 536
rect -2241 487 -2229 521
rect -2195 487 -2183 521
rect -2241 453 -2183 487
rect -2241 419 -2229 453
rect -2195 419 -2183 453
rect -2241 385 -2183 419
rect -2241 351 -2229 385
rect -2195 351 -2183 385
rect -2241 336 -2183 351
rect -2083 521 -2025 536
rect -2083 487 -2071 521
rect -2037 487 -2025 521
rect -2083 453 -2025 487
rect -2083 419 -2071 453
rect -2037 419 -2025 453
rect -2083 385 -2025 419
rect -2083 351 -2071 385
rect -2037 351 -2025 385
rect -2083 336 -2025 351
rect -1925 521 -1867 536
rect -1925 487 -1913 521
rect -1879 487 -1867 521
rect -1925 453 -1867 487
rect -1925 419 -1913 453
rect -1879 419 -1867 453
rect -1925 385 -1867 419
rect -1925 351 -1913 385
rect -1879 351 -1867 385
rect -1925 336 -1867 351
rect -1767 521 -1709 536
rect -1767 487 -1755 521
rect -1721 487 -1709 521
rect -1767 453 -1709 487
rect -1767 419 -1755 453
rect -1721 419 -1709 453
rect -1767 385 -1709 419
rect -1767 351 -1755 385
rect -1721 351 -1709 385
rect -1767 336 -1709 351
rect -1609 521 -1551 536
rect -1609 487 -1597 521
rect -1563 487 -1551 521
rect -1609 453 -1551 487
rect -1609 419 -1597 453
rect -1563 419 -1551 453
rect -1609 385 -1551 419
rect -1609 351 -1597 385
rect -1563 351 -1551 385
rect -1609 336 -1551 351
rect -1451 521 -1393 536
rect -1451 487 -1439 521
rect -1405 487 -1393 521
rect -1451 453 -1393 487
rect -1451 419 -1439 453
rect -1405 419 -1393 453
rect -1451 385 -1393 419
rect -1451 351 -1439 385
rect -1405 351 -1393 385
rect -1451 336 -1393 351
rect -1293 521 -1235 536
rect -1293 487 -1281 521
rect -1247 487 -1235 521
rect -1293 453 -1235 487
rect -1293 419 -1281 453
rect -1247 419 -1235 453
rect -1293 385 -1235 419
rect -1293 351 -1281 385
rect -1247 351 -1235 385
rect -1293 336 -1235 351
rect -1135 521 -1077 536
rect -1135 487 -1123 521
rect -1089 487 -1077 521
rect -1135 453 -1077 487
rect -1135 419 -1123 453
rect -1089 419 -1077 453
rect -1135 385 -1077 419
rect -1135 351 -1123 385
rect -1089 351 -1077 385
rect -1135 336 -1077 351
rect -977 521 -919 536
rect -977 487 -965 521
rect -931 487 -919 521
rect -977 453 -919 487
rect -977 419 -965 453
rect -931 419 -919 453
rect -977 385 -919 419
rect -977 351 -965 385
rect -931 351 -919 385
rect -977 336 -919 351
rect -819 521 -761 536
rect -819 487 -807 521
rect -773 487 -761 521
rect -819 453 -761 487
rect -819 419 -807 453
rect -773 419 -761 453
rect -819 385 -761 419
rect -819 351 -807 385
rect -773 351 -761 385
rect -819 336 -761 351
rect -661 521 -603 536
rect -661 487 -649 521
rect -615 487 -603 521
rect -661 453 -603 487
rect -661 419 -649 453
rect -615 419 -603 453
rect -661 385 -603 419
rect -661 351 -649 385
rect -615 351 -603 385
rect -661 336 -603 351
rect -503 521 -445 536
rect -503 487 -491 521
rect -457 487 -445 521
rect -503 453 -445 487
rect -503 419 -491 453
rect -457 419 -445 453
rect -503 385 -445 419
rect -503 351 -491 385
rect -457 351 -445 385
rect -503 336 -445 351
rect -345 521 -287 536
rect -345 487 -333 521
rect -299 487 -287 521
rect -345 453 -287 487
rect -345 419 -333 453
rect -299 419 -287 453
rect -345 385 -287 419
rect -345 351 -333 385
rect -299 351 -287 385
rect -345 336 -287 351
rect -187 521 -129 536
rect -187 487 -175 521
rect -141 487 -129 521
rect -187 453 -129 487
rect -187 419 -175 453
rect -141 419 -129 453
rect -187 385 -129 419
rect -187 351 -175 385
rect -141 351 -129 385
rect -187 336 -129 351
rect -29 521 29 536
rect -29 487 -17 521
rect 17 487 29 521
rect -29 453 29 487
rect -29 419 -17 453
rect 17 419 29 453
rect -29 385 29 419
rect -29 351 -17 385
rect 17 351 29 385
rect -29 336 29 351
rect 129 521 187 536
rect 129 487 141 521
rect 175 487 187 521
rect 129 453 187 487
rect 129 419 141 453
rect 175 419 187 453
rect 129 385 187 419
rect 129 351 141 385
rect 175 351 187 385
rect 129 336 187 351
rect 287 521 345 536
rect 287 487 299 521
rect 333 487 345 521
rect 287 453 345 487
rect 287 419 299 453
rect 333 419 345 453
rect 287 385 345 419
rect 287 351 299 385
rect 333 351 345 385
rect 287 336 345 351
rect 445 521 503 536
rect 445 487 457 521
rect 491 487 503 521
rect 445 453 503 487
rect 445 419 457 453
rect 491 419 503 453
rect 445 385 503 419
rect 445 351 457 385
rect 491 351 503 385
rect 445 336 503 351
rect 603 521 661 536
rect 603 487 615 521
rect 649 487 661 521
rect 603 453 661 487
rect 603 419 615 453
rect 649 419 661 453
rect 603 385 661 419
rect 603 351 615 385
rect 649 351 661 385
rect 603 336 661 351
rect 761 521 819 536
rect 761 487 773 521
rect 807 487 819 521
rect 761 453 819 487
rect 761 419 773 453
rect 807 419 819 453
rect 761 385 819 419
rect 761 351 773 385
rect 807 351 819 385
rect 761 336 819 351
rect 919 521 977 536
rect 919 487 931 521
rect 965 487 977 521
rect 919 453 977 487
rect 919 419 931 453
rect 965 419 977 453
rect 919 385 977 419
rect 919 351 931 385
rect 965 351 977 385
rect 919 336 977 351
rect 1077 521 1135 536
rect 1077 487 1089 521
rect 1123 487 1135 521
rect 1077 453 1135 487
rect 1077 419 1089 453
rect 1123 419 1135 453
rect 1077 385 1135 419
rect 1077 351 1089 385
rect 1123 351 1135 385
rect 1077 336 1135 351
rect 1235 521 1293 536
rect 1235 487 1247 521
rect 1281 487 1293 521
rect 1235 453 1293 487
rect 1235 419 1247 453
rect 1281 419 1293 453
rect 1235 385 1293 419
rect 1235 351 1247 385
rect 1281 351 1293 385
rect 1235 336 1293 351
rect 1393 521 1451 536
rect 1393 487 1405 521
rect 1439 487 1451 521
rect 1393 453 1451 487
rect 1393 419 1405 453
rect 1439 419 1451 453
rect 1393 385 1451 419
rect 1393 351 1405 385
rect 1439 351 1451 385
rect 1393 336 1451 351
rect 1551 521 1609 536
rect 1551 487 1563 521
rect 1597 487 1609 521
rect 1551 453 1609 487
rect 1551 419 1563 453
rect 1597 419 1609 453
rect 1551 385 1609 419
rect 1551 351 1563 385
rect 1597 351 1609 385
rect 1551 336 1609 351
rect 1709 521 1767 536
rect 1709 487 1721 521
rect 1755 487 1767 521
rect 1709 453 1767 487
rect 1709 419 1721 453
rect 1755 419 1767 453
rect 1709 385 1767 419
rect 1709 351 1721 385
rect 1755 351 1767 385
rect 1709 336 1767 351
rect 1867 521 1925 536
rect 1867 487 1879 521
rect 1913 487 1925 521
rect 1867 453 1925 487
rect 1867 419 1879 453
rect 1913 419 1925 453
rect 1867 385 1925 419
rect 1867 351 1879 385
rect 1913 351 1925 385
rect 1867 336 1925 351
rect 2025 521 2083 536
rect 2025 487 2037 521
rect 2071 487 2083 521
rect 2025 453 2083 487
rect 2025 419 2037 453
rect 2071 419 2083 453
rect 2025 385 2083 419
rect 2025 351 2037 385
rect 2071 351 2083 385
rect 2025 336 2083 351
rect 2183 521 2241 536
rect 2183 487 2195 521
rect 2229 487 2241 521
rect 2183 453 2241 487
rect 2183 419 2195 453
rect 2229 419 2241 453
rect 2183 385 2241 419
rect 2183 351 2195 385
rect 2229 351 2241 385
rect 2183 336 2241 351
rect 2341 521 2399 536
rect 2341 487 2353 521
rect 2387 487 2399 521
rect 2341 453 2399 487
rect 2341 419 2353 453
rect 2387 419 2399 453
rect 2341 385 2399 419
rect 2341 351 2353 385
rect 2387 351 2399 385
rect 2341 336 2399 351
rect 2499 521 2557 536
rect 2499 487 2511 521
rect 2545 487 2557 521
rect 2499 453 2557 487
rect 2499 419 2511 453
rect 2545 419 2557 453
rect 2499 385 2557 419
rect 2499 351 2511 385
rect 2545 351 2557 385
rect 2499 336 2557 351
rect 2657 521 2715 536
rect 2657 487 2669 521
rect 2703 487 2715 521
rect 2657 453 2715 487
rect 2657 419 2669 453
rect 2703 419 2715 453
rect 2657 385 2715 419
rect 2657 351 2669 385
rect 2703 351 2715 385
rect 2657 336 2715 351
rect 2815 521 2873 536
rect 2815 487 2827 521
rect 2861 487 2873 521
rect 2815 453 2873 487
rect 2815 419 2827 453
rect 2861 419 2873 453
rect 2815 385 2873 419
rect 2815 351 2827 385
rect 2861 351 2873 385
rect 2815 336 2873 351
rect 2973 521 3031 536
rect 2973 487 2985 521
rect 3019 487 3031 521
rect 2973 453 3031 487
rect 2973 419 2985 453
rect 3019 419 3031 453
rect 2973 385 3031 419
rect 2973 351 2985 385
rect 3019 351 3031 385
rect 2973 336 3031 351
rect 3131 521 3189 536
rect 3131 487 3143 521
rect 3177 487 3189 521
rect 3131 453 3189 487
rect 3131 419 3143 453
rect 3177 419 3189 453
rect 3131 385 3189 419
rect 3131 351 3143 385
rect 3177 351 3189 385
rect 3131 336 3189 351
rect -3189 85 -3131 100
rect -3189 51 -3177 85
rect -3143 51 -3131 85
rect -3189 17 -3131 51
rect -3189 -17 -3177 17
rect -3143 -17 -3131 17
rect -3189 -51 -3131 -17
rect -3189 -85 -3177 -51
rect -3143 -85 -3131 -51
rect -3189 -100 -3131 -85
rect -3031 85 -2973 100
rect -3031 51 -3019 85
rect -2985 51 -2973 85
rect -3031 17 -2973 51
rect -3031 -17 -3019 17
rect -2985 -17 -2973 17
rect -3031 -51 -2973 -17
rect -3031 -85 -3019 -51
rect -2985 -85 -2973 -51
rect -3031 -100 -2973 -85
rect -2873 85 -2815 100
rect -2873 51 -2861 85
rect -2827 51 -2815 85
rect -2873 17 -2815 51
rect -2873 -17 -2861 17
rect -2827 -17 -2815 17
rect -2873 -51 -2815 -17
rect -2873 -85 -2861 -51
rect -2827 -85 -2815 -51
rect -2873 -100 -2815 -85
rect -2715 85 -2657 100
rect -2715 51 -2703 85
rect -2669 51 -2657 85
rect -2715 17 -2657 51
rect -2715 -17 -2703 17
rect -2669 -17 -2657 17
rect -2715 -51 -2657 -17
rect -2715 -85 -2703 -51
rect -2669 -85 -2657 -51
rect -2715 -100 -2657 -85
rect -2557 85 -2499 100
rect -2557 51 -2545 85
rect -2511 51 -2499 85
rect -2557 17 -2499 51
rect -2557 -17 -2545 17
rect -2511 -17 -2499 17
rect -2557 -51 -2499 -17
rect -2557 -85 -2545 -51
rect -2511 -85 -2499 -51
rect -2557 -100 -2499 -85
rect -2399 85 -2341 100
rect -2399 51 -2387 85
rect -2353 51 -2341 85
rect -2399 17 -2341 51
rect -2399 -17 -2387 17
rect -2353 -17 -2341 17
rect -2399 -51 -2341 -17
rect -2399 -85 -2387 -51
rect -2353 -85 -2341 -51
rect -2399 -100 -2341 -85
rect -2241 85 -2183 100
rect -2241 51 -2229 85
rect -2195 51 -2183 85
rect -2241 17 -2183 51
rect -2241 -17 -2229 17
rect -2195 -17 -2183 17
rect -2241 -51 -2183 -17
rect -2241 -85 -2229 -51
rect -2195 -85 -2183 -51
rect -2241 -100 -2183 -85
rect -2083 85 -2025 100
rect -2083 51 -2071 85
rect -2037 51 -2025 85
rect -2083 17 -2025 51
rect -2083 -17 -2071 17
rect -2037 -17 -2025 17
rect -2083 -51 -2025 -17
rect -2083 -85 -2071 -51
rect -2037 -85 -2025 -51
rect -2083 -100 -2025 -85
rect -1925 85 -1867 100
rect -1925 51 -1913 85
rect -1879 51 -1867 85
rect -1925 17 -1867 51
rect -1925 -17 -1913 17
rect -1879 -17 -1867 17
rect -1925 -51 -1867 -17
rect -1925 -85 -1913 -51
rect -1879 -85 -1867 -51
rect -1925 -100 -1867 -85
rect -1767 85 -1709 100
rect -1767 51 -1755 85
rect -1721 51 -1709 85
rect -1767 17 -1709 51
rect -1767 -17 -1755 17
rect -1721 -17 -1709 17
rect -1767 -51 -1709 -17
rect -1767 -85 -1755 -51
rect -1721 -85 -1709 -51
rect -1767 -100 -1709 -85
rect -1609 85 -1551 100
rect -1609 51 -1597 85
rect -1563 51 -1551 85
rect -1609 17 -1551 51
rect -1609 -17 -1597 17
rect -1563 -17 -1551 17
rect -1609 -51 -1551 -17
rect -1609 -85 -1597 -51
rect -1563 -85 -1551 -51
rect -1609 -100 -1551 -85
rect -1451 85 -1393 100
rect -1451 51 -1439 85
rect -1405 51 -1393 85
rect -1451 17 -1393 51
rect -1451 -17 -1439 17
rect -1405 -17 -1393 17
rect -1451 -51 -1393 -17
rect -1451 -85 -1439 -51
rect -1405 -85 -1393 -51
rect -1451 -100 -1393 -85
rect -1293 85 -1235 100
rect -1293 51 -1281 85
rect -1247 51 -1235 85
rect -1293 17 -1235 51
rect -1293 -17 -1281 17
rect -1247 -17 -1235 17
rect -1293 -51 -1235 -17
rect -1293 -85 -1281 -51
rect -1247 -85 -1235 -51
rect -1293 -100 -1235 -85
rect -1135 85 -1077 100
rect -1135 51 -1123 85
rect -1089 51 -1077 85
rect -1135 17 -1077 51
rect -1135 -17 -1123 17
rect -1089 -17 -1077 17
rect -1135 -51 -1077 -17
rect -1135 -85 -1123 -51
rect -1089 -85 -1077 -51
rect -1135 -100 -1077 -85
rect -977 85 -919 100
rect -977 51 -965 85
rect -931 51 -919 85
rect -977 17 -919 51
rect -977 -17 -965 17
rect -931 -17 -919 17
rect -977 -51 -919 -17
rect -977 -85 -965 -51
rect -931 -85 -919 -51
rect -977 -100 -919 -85
rect -819 85 -761 100
rect -819 51 -807 85
rect -773 51 -761 85
rect -819 17 -761 51
rect -819 -17 -807 17
rect -773 -17 -761 17
rect -819 -51 -761 -17
rect -819 -85 -807 -51
rect -773 -85 -761 -51
rect -819 -100 -761 -85
rect -661 85 -603 100
rect -661 51 -649 85
rect -615 51 -603 85
rect -661 17 -603 51
rect -661 -17 -649 17
rect -615 -17 -603 17
rect -661 -51 -603 -17
rect -661 -85 -649 -51
rect -615 -85 -603 -51
rect -661 -100 -603 -85
rect -503 85 -445 100
rect -503 51 -491 85
rect -457 51 -445 85
rect -503 17 -445 51
rect -503 -17 -491 17
rect -457 -17 -445 17
rect -503 -51 -445 -17
rect -503 -85 -491 -51
rect -457 -85 -445 -51
rect -503 -100 -445 -85
rect -345 85 -287 100
rect -345 51 -333 85
rect -299 51 -287 85
rect -345 17 -287 51
rect -345 -17 -333 17
rect -299 -17 -287 17
rect -345 -51 -287 -17
rect -345 -85 -333 -51
rect -299 -85 -287 -51
rect -345 -100 -287 -85
rect -187 85 -129 100
rect -187 51 -175 85
rect -141 51 -129 85
rect -187 17 -129 51
rect -187 -17 -175 17
rect -141 -17 -129 17
rect -187 -51 -129 -17
rect -187 -85 -175 -51
rect -141 -85 -129 -51
rect -187 -100 -129 -85
rect -29 85 29 100
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -100 29 -85
rect 129 85 187 100
rect 129 51 141 85
rect 175 51 187 85
rect 129 17 187 51
rect 129 -17 141 17
rect 175 -17 187 17
rect 129 -51 187 -17
rect 129 -85 141 -51
rect 175 -85 187 -51
rect 129 -100 187 -85
rect 287 85 345 100
rect 287 51 299 85
rect 333 51 345 85
rect 287 17 345 51
rect 287 -17 299 17
rect 333 -17 345 17
rect 287 -51 345 -17
rect 287 -85 299 -51
rect 333 -85 345 -51
rect 287 -100 345 -85
rect 445 85 503 100
rect 445 51 457 85
rect 491 51 503 85
rect 445 17 503 51
rect 445 -17 457 17
rect 491 -17 503 17
rect 445 -51 503 -17
rect 445 -85 457 -51
rect 491 -85 503 -51
rect 445 -100 503 -85
rect 603 85 661 100
rect 603 51 615 85
rect 649 51 661 85
rect 603 17 661 51
rect 603 -17 615 17
rect 649 -17 661 17
rect 603 -51 661 -17
rect 603 -85 615 -51
rect 649 -85 661 -51
rect 603 -100 661 -85
rect 761 85 819 100
rect 761 51 773 85
rect 807 51 819 85
rect 761 17 819 51
rect 761 -17 773 17
rect 807 -17 819 17
rect 761 -51 819 -17
rect 761 -85 773 -51
rect 807 -85 819 -51
rect 761 -100 819 -85
rect 919 85 977 100
rect 919 51 931 85
rect 965 51 977 85
rect 919 17 977 51
rect 919 -17 931 17
rect 965 -17 977 17
rect 919 -51 977 -17
rect 919 -85 931 -51
rect 965 -85 977 -51
rect 919 -100 977 -85
rect 1077 85 1135 100
rect 1077 51 1089 85
rect 1123 51 1135 85
rect 1077 17 1135 51
rect 1077 -17 1089 17
rect 1123 -17 1135 17
rect 1077 -51 1135 -17
rect 1077 -85 1089 -51
rect 1123 -85 1135 -51
rect 1077 -100 1135 -85
rect 1235 85 1293 100
rect 1235 51 1247 85
rect 1281 51 1293 85
rect 1235 17 1293 51
rect 1235 -17 1247 17
rect 1281 -17 1293 17
rect 1235 -51 1293 -17
rect 1235 -85 1247 -51
rect 1281 -85 1293 -51
rect 1235 -100 1293 -85
rect 1393 85 1451 100
rect 1393 51 1405 85
rect 1439 51 1451 85
rect 1393 17 1451 51
rect 1393 -17 1405 17
rect 1439 -17 1451 17
rect 1393 -51 1451 -17
rect 1393 -85 1405 -51
rect 1439 -85 1451 -51
rect 1393 -100 1451 -85
rect 1551 85 1609 100
rect 1551 51 1563 85
rect 1597 51 1609 85
rect 1551 17 1609 51
rect 1551 -17 1563 17
rect 1597 -17 1609 17
rect 1551 -51 1609 -17
rect 1551 -85 1563 -51
rect 1597 -85 1609 -51
rect 1551 -100 1609 -85
rect 1709 85 1767 100
rect 1709 51 1721 85
rect 1755 51 1767 85
rect 1709 17 1767 51
rect 1709 -17 1721 17
rect 1755 -17 1767 17
rect 1709 -51 1767 -17
rect 1709 -85 1721 -51
rect 1755 -85 1767 -51
rect 1709 -100 1767 -85
rect 1867 85 1925 100
rect 1867 51 1879 85
rect 1913 51 1925 85
rect 1867 17 1925 51
rect 1867 -17 1879 17
rect 1913 -17 1925 17
rect 1867 -51 1925 -17
rect 1867 -85 1879 -51
rect 1913 -85 1925 -51
rect 1867 -100 1925 -85
rect 2025 85 2083 100
rect 2025 51 2037 85
rect 2071 51 2083 85
rect 2025 17 2083 51
rect 2025 -17 2037 17
rect 2071 -17 2083 17
rect 2025 -51 2083 -17
rect 2025 -85 2037 -51
rect 2071 -85 2083 -51
rect 2025 -100 2083 -85
rect 2183 85 2241 100
rect 2183 51 2195 85
rect 2229 51 2241 85
rect 2183 17 2241 51
rect 2183 -17 2195 17
rect 2229 -17 2241 17
rect 2183 -51 2241 -17
rect 2183 -85 2195 -51
rect 2229 -85 2241 -51
rect 2183 -100 2241 -85
rect 2341 85 2399 100
rect 2341 51 2353 85
rect 2387 51 2399 85
rect 2341 17 2399 51
rect 2341 -17 2353 17
rect 2387 -17 2399 17
rect 2341 -51 2399 -17
rect 2341 -85 2353 -51
rect 2387 -85 2399 -51
rect 2341 -100 2399 -85
rect 2499 85 2557 100
rect 2499 51 2511 85
rect 2545 51 2557 85
rect 2499 17 2557 51
rect 2499 -17 2511 17
rect 2545 -17 2557 17
rect 2499 -51 2557 -17
rect 2499 -85 2511 -51
rect 2545 -85 2557 -51
rect 2499 -100 2557 -85
rect 2657 85 2715 100
rect 2657 51 2669 85
rect 2703 51 2715 85
rect 2657 17 2715 51
rect 2657 -17 2669 17
rect 2703 -17 2715 17
rect 2657 -51 2715 -17
rect 2657 -85 2669 -51
rect 2703 -85 2715 -51
rect 2657 -100 2715 -85
rect 2815 85 2873 100
rect 2815 51 2827 85
rect 2861 51 2873 85
rect 2815 17 2873 51
rect 2815 -17 2827 17
rect 2861 -17 2873 17
rect 2815 -51 2873 -17
rect 2815 -85 2827 -51
rect 2861 -85 2873 -51
rect 2815 -100 2873 -85
rect 2973 85 3031 100
rect 2973 51 2985 85
rect 3019 51 3031 85
rect 2973 17 3031 51
rect 2973 -17 2985 17
rect 3019 -17 3031 17
rect 2973 -51 3031 -17
rect 2973 -85 2985 -51
rect 3019 -85 3031 -51
rect 2973 -100 3031 -85
rect 3131 85 3189 100
rect 3131 51 3143 85
rect 3177 51 3189 85
rect 3131 17 3189 51
rect 3131 -17 3143 17
rect 3177 -17 3189 17
rect 3131 -51 3189 -17
rect 3131 -85 3143 -51
rect 3177 -85 3189 -51
rect 3131 -100 3189 -85
rect -3189 -351 -3131 -336
rect -3189 -385 -3177 -351
rect -3143 -385 -3131 -351
rect -3189 -419 -3131 -385
rect -3189 -453 -3177 -419
rect -3143 -453 -3131 -419
rect -3189 -487 -3131 -453
rect -3189 -521 -3177 -487
rect -3143 -521 -3131 -487
rect -3189 -536 -3131 -521
rect -3031 -351 -2973 -336
rect -3031 -385 -3019 -351
rect -2985 -385 -2973 -351
rect -3031 -419 -2973 -385
rect -3031 -453 -3019 -419
rect -2985 -453 -2973 -419
rect -3031 -487 -2973 -453
rect -3031 -521 -3019 -487
rect -2985 -521 -2973 -487
rect -3031 -536 -2973 -521
rect -2873 -351 -2815 -336
rect -2873 -385 -2861 -351
rect -2827 -385 -2815 -351
rect -2873 -419 -2815 -385
rect -2873 -453 -2861 -419
rect -2827 -453 -2815 -419
rect -2873 -487 -2815 -453
rect -2873 -521 -2861 -487
rect -2827 -521 -2815 -487
rect -2873 -536 -2815 -521
rect -2715 -351 -2657 -336
rect -2715 -385 -2703 -351
rect -2669 -385 -2657 -351
rect -2715 -419 -2657 -385
rect -2715 -453 -2703 -419
rect -2669 -453 -2657 -419
rect -2715 -487 -2657 -453
rect -2715 -521 -2703 -487
rect -2669 -521 -2657 -487
rect -2715 -536 -2657 -521
rect -2557 -351 -2499 -336
rect -2557 -385 -2545 -351
rect -2511 -385 -2499 -351
rect -2557 -419 -2499 -385
rect -2557 -453 -2545 -419
rect -2511 -453 -2499 -419
rect -2557 -487 -2499 -453
rect -2557 -521 -2545 -487
rect -2511 -521 -2499 -487
rect -2557 -536 -2499 -521
rect -2399 -351 -2341 -336
rect -2399 -385 -2387 -351
rect -2353 -385 -2341 -351
rect -2399 -419 -2341 -385
rect -2399 -453 -2387 -419
rect -2353 -453 -2341 -419
rect -2399 -487 -2341 -453
rect -2399 -521 -2387 -487
rect -2353 -521 -2341 -487
rect -2399 -536 -2341 -521
rect -2241 -351 -2183 -336
rect -2241 -385 -2229 -351
rect -2195 -385 -2183 -351
rect -2241 -419 -2183 -385
rect -2241 -453 -2229 -419
rect -2195 -453 -2183 -419
rect -2241 -487 -2183 -453
rect -2241 -521 -2229 -487
rect -2195 -521 -2183 -487
rect -2241 -536 -2183 -521
rect -2083 -351 -2025 -336
rect -2083 -385 -2071 -351
rect -2037 -385 -2025 -351
rect -2083 -419 -2025 -385
rect -2083 -453 -2071 -419
rect -2037 -453 -2025 -419
rect -2083 -487 -2025 -453
rect -2083 -521 -2071 -487
rect -2037 -521 -2025 -487
rect -2083 -536 -2025 -521
rect -1925 -351 -1867 -336
rect -1925 -385 -1913 -351
rect -1879 -385 -1867 -351
rect -1925 -419 -1867 -385
rect -1925 -453 -1913 -419
rect -1879 -453 -1867 -419
rect -1925 -487 -1867 -453
rect -1925 -521 -1913 -487
rect -1879 -521 -1867 -487
rect -1925 -536 -1867 -521
rect -1767 -351 -1709 -336
rect -1767 -385 -1755 -351
rect -1721 -385 -1709 -351
rect -1767 -419 -1709 -385
rect -1767 -453 -1755 -419
rect -1721 -453 -1709 -419
rect -1767 -487 -1709 -453
rect -1767 -521 -1755 -487
rect -1721 -521 -1709 -487
rect -1767 -536 -1709 -521
rect -1609 -351 -1551 -336
rect -1609 -385 -1597 -351
rect -1563 -385 -1551 -351
rect -1609 -419 -1551 -385
rect -1609 -453 -1597 -419
rect -1563 -453 -1551 -419
rect -1609 -487 -1551 -453
rect -1609 -521 -1597 -487
rect -1563 -521 -1551 -487
rect -1609 -536 -1551 -521
rect -1451 -351 -1393 -336
rect -1451 -385 -1439 -351
rect -1405 -385 -1393 -351
rect -1451 -419 -1393 -385
rect -1451 -453 -1439 -419
rect -1405 -453 -1393 -419
rect -1451 -487 -1393 -453
rect -1451 -521 -1439 -487
rect -1405 -521 -1393 -487
rect -1451 -536 -1393 -521
rect -1293 -351 -1235 -336
rect -1293 -385 -1281 -351
rect -1247 -385 -1235 -351
rect -1293 -419 -1235 -385
rect -1293 -453 -1281 -419
rect -1247 -453 -1235 -419
rect -1293 -487 -1235 -453
rect -1293 -521 -1281 -487
rect -1247 -521 -1235 -487
rect -1293 -536 -1235 -521
rect -1135 -351 -1077 -336
rect -1135 -385 -1123 -351
rect -1089 -385 -1077 -351
rect -1135 -419 -1077 -385
rect -1135 -453 -1123 -419
rect -1089 -453 -1077 -419
rect -1135 -487 -1077 -453
rect -1135 -521 -1123 -487
rect -1089 -521 -1077 -487
rect -1135 -536 -1077 -521
rect -977 -351 -919 -336
rect -977 -385 -965 -351
rect -931 -385 -919 -351
rect -977 -419 -919 -385
rect -977 -453 -965 -419
rect -931 -453 -919 -419
rect -977 -487 -919 -453
rect -977 -521 -965 -487
rect -931 -521 -919 -487
rect -977 -536 -919 -521
rect -819 -351 -761 -336
rect -819 -385 -807 -351
rect -773 -385 -761 -351
rect -819 -419 -761 -385
rect -819 -453 -807 -419
rect -773 -453 -761 -419
rect -819 -487 -761 -453
rect -819 -521 -807 -487
rect -773 -521 -761 -487
rect -819 -536 -761 -521
rect -661 -351 -603 -336
rect -661 -385 -649 -351
rect -615 -385 -603 -351
rect -661 -419 -603 -385
rect -661 -453 -649 -419
rect -615 -453 -603 -419
rect -661 -487 -603 -453
rect -661 -521 -649 -487
rect -615 -521 -603 -487
rect -661 -536 -603 -521
rect -503 -351 -445 -336
rect -503 -385 -491 -351
rect -457 -385 -445 -351
rect -503 -419 -445 -385
rect -503 -453 -491 -419
rect -457 -453 -445 -419
rect -503 -487 -445 -453
rect -503 -521 -491 -487
rect -457 -521 -445 -487
rect -503 -536 -445 -521
rect -345 -351 -287 -336
rect -345 -385 -333 -351
rect -299 -385 -287 -351
rect -345 -419 -287 -385
rect -345 -453 -333 -419
rect -299 -453 -287 -419
rect -345 -487 -287 -453
rect -345 -521 -333 -487
rect -299 -521 -287 -487
rect -345 -536 -287 -521
rect -187 -351 -129 -336
rect -187 -385 -175 -351
rect -141 -385 -129 -351
rect -187 -419 -129 -385
rect -187 -453 -175 -419
rect -141 -453 -129 -419
rect -187 -487 -129 -453
rect -187 -521 -175 -487
rect -141 -521 -129 -487
rect -187 -536 -129 -521
rect -29 -351 29 -336
rect -29 -385 -17 -351
rect 17 -385 29 -351
rect -29 -419 29 -385
rect -29 -453 -17 -419
rect 17 -453 29 -419
rect -29 -487 29 -453
rect -29 -521 -17 -487
rect 17 -521 29 -487
rect -29 -536 29 -521
rect 129 -351 187 -336
rect 129 -385 141 -351
rect 175 -385 187 -351
rect 129 -419 187 -385
rect 129 -453 141 -419
rect 175 -453 187 -419
rect 129 -487 187 -453
rect 129 -521 141 -487
rect 175 -521 187 -487
rect 129 -536 187 -521
rect 287 -351 345 -336
rect 287 -385 299 -351
rect 333 -385 345 -351
rect 287 -419 345 -385
rect 287 -453 299 -419
rect 333 -453 345 -419
rect 287 -487 345 -453
rect 287 -521 299 -487
rect 333 -521 345 -487
rect 287 -536 345 -521
rect 445 -351 503 -336
rect 445 -385 457 -351
rect 491 -385 503 -351
rect 445 -419 503 -385
rect 445 -453 457 -419
rect 491 -453 503 -419
rect 445 -487 503 -453
rect 445 -521 457 -487
rect 491 -521 503 -487
rect 445 -536 503 -521
rect 603 -351 661 -336
rect 603 -385 615 -351
rect 649 -385 661 -351
rect 603 -419 661 -385
rect 603 -453 615 -419
rect 649 -453 661 -419
rect 603 -487 661 -453
rect 603 -521 615 -487
rect 649 -521 661 -487
rect 603 -536 661 -521
rect 761 -351 819 -336
rect 761 -385 773 -351
rect 807 -385 819 -351
rect 761 -419 819 -385
rect 761 -453 773 -419
rect 807 -453 819 -419
rect 761 -487 819 -453
rect 761 -521 773 -487
rect 807 -521 819 -487
rect 761 -536 819 -521
rect 919 -351 977 -336
rect 919 -385 931 -351
rect 965 -385 977 -351
rect 919 -419 977 -385
rect 919 -453 931 -419
rect 965 -453 977 -419
rect 919 -487 977 -453
rect 919 -521 931 -487
rect 965 -521 977 -487
rect 919 -536 977 -521
rect 1077 -351 1135 -336
rect 1077 -385 1089 -351
rect 1123 -385 1135 -351
rect 1077 -419 1135 -385
rect 1077 -453 1089 -419
rect 1123 -453 1135 -419
rect 1077 -487 1135 -453
rect 1077 -521 1089 -487
rect 1123 -521 1135 -487
rect 1077 -536 1135 -521
rect 1235 -351 1293 -336
rect 1235 -385 1247 -351
rect 1281 -385 1293 -351
rect 1235 -419 1293 -385
rect 1235 -453 1247 -419
rect 1281 -453 1293 -419
rect 1235 -487 1293 -453
rect 1235 -521 1247 -487
rect 1281 -521 1293 -487
rect 1235 -536 1293 -521
rect 1393 -351 1451 -336
rect 1393 -385 1405 -351
rect 1439 -385 1451 -351
rect 1393 -419 1451 -385
rect 1393 -453 1405 -419
rect 1439 -453 1451 -419
rect 1393 -487 1451 -453
rect 1393 -521 1405 -487
rect 1439 -521 1451 -487
rect 1393 -536 1451 -521
rect 1551 -351 1609 -336
rect 1551 -385 1563 -351
rect 1597 -385 1609 -351
rect 1551 -419 1609 -385
rect 1551 -453 1563 -419
rect 1597 -453 1609 -419
rect 1551 -487 1609 -453
rect 1551 -521 1563 -487
rect 1597 -521 1609 -487
rect 1551 -536 1609 -521
rect 1709 -351 1767 -336
rect 1709 -385 1721 -351
rect 1755 -385 1767 -351
rect 1709 -419 1767 -385
rect 1709 -453 1721 -419
rect 1755 -453 1767 -419
rect 1709 -487 1767 -453
rect 1709 -521 1721 -487
rect 1755 -521 1767 -487
rect 1709 -536 1767 -521
rect 1867 -351 1925 -336
rect 1867 -385 1879 -351
rect 1913 -385 1925 -351
rect 1867 -419 1925 -385
rect 1867 -453 1879 -419
rect 1913 -453 1925 -419
rect 1867 -487 1925 -453
rect 1867 -521 1879 -487
rect 1913 -521 1925 -487
rect 1867 -536 1925 -521
rect 2025 -351 2083 -336
rect 2025 -385 2037 -351
rect 2071 -385 2083 -351
rect 2025 -419 2083 -385
rect 2025 -453 2037 -419
rect 2071 -453 2083 -419
rect 2025 -487 2083 -453
rect 2025 -521 2037 -487
rect 2071 -521 2083 -487
rect 2025 -536 2083 -521
rect 2183 -351 2241 -336
rect 2183 -385 2195 -351
rect 2229 -385 2241 -351
rect 2183 -419 2241 -385
rect 2183 -453 2195 -419
rect 2229 -453 2241 -419
rect 2183 -487 2241 -453
rect 2183 -521 2195 -487
rect 2229 -521 2241 -487
rect 2183 -536 2241 -521
rect 2341 -351 2399 -336
rect 2341 -385 2353 -351
rect 2387 -385 2399 -351
rect 2341 -419 2399 -385
rect 2341 -453 2353 -419
rect 2387 -453 2399 -419
rect 2341 -487 2399 -453
rect 2341 -521 2353 -487
rect 2387 -521 2399 -487
rect 2341 -536 2399 -521
rect 2499 -351 2557 -336
rect 2499 -385 2511 -351
rect 2545 -385 2557 -351
rect 2499 -419 2557 -385
rect 2499 -453 2511 -419
rect 2545 -453 2557 -419
rect 2499 -487 2557 -453
rect 2499 -521 2511 -487
rect 2545 -521 2557 -487
rect 2499 -536 2557 -521
rect 2657 -351 2715 -336
rect 2657 -385 2669 -351
rect 2703 -385 2715 -351
rect 2657 -419 2715 -385
rect 2657 -453 2669 -419
rect 2703 -453 2715 -419
rect 2657 -487 2715 -453
rect 2657 -521 2669 -487
rect 2703 -521 2715 -487
rect 2657 -536 2715 -521
rect 2815 -351 2873 -336
rect 2815 -385 2827 -351
rect 2861 -385 2873 -351
rect 2815 -419 2873 -385
rect 2815 -453 2827 -419
rect 2861 -453 2873 -419
rect 2815 -487 2873 -453
rect 2815 -521 2827 -487
rect 2861 -521 2873 -487
rect 2815 -536 2873 -521
rect 2973 -351 3031 -336
rect 2973 -385 2985 -351
rect 3019 -385 3031 -351
rect 2973 -419 3031 -385
rect 2973 -453 2985 -419
rect 3019 -453 3031 -419
rect 2973 -487 3031 -453
rect 2973 -521 2985 -487
rect 3019 -521 3031 -487
rect 2973 -536 3031 -521
rect 3131 -351 3189 -336
rect 3131 -385 3143 -351
rect 3177 -385 3189 -351
rect 3131 -419 3189 -385
rect 3131 -453 3143 -419
rect 3177 -453 3189 -419
rect 3131 -487 3189 -453
rect 3131 -521 3143 -487
rect 3177 -521 3189 -487
rect 3131 -536 3189 -521
rect -3189 -787 -3131 -772
rect -3189 -821 -3177 -787
rect -3143 -821 -3131 -787
rect -3189 -855 -3131 -821
rect -3189 -889 -3177 -855
rect -3143 -889 -3131 -855
rect -3189 -923 -3131 -889
rect -3189 -957 -3177 -923
rect -3143 -957 -3131 -923
rect -3189 -972 -3131 -957
rect -3031 -787 -2973 -772
rect -3031 -821 -3019 -787
rect -2985 -821 -2973 -787
rect -3031 -855 -2973 -821
rect -3031 -889 -3019 -855
rect -2985 -889 -2973 -855
rect -3031 -923 -2973 -889
rect -3031 -957 -3019 -923
rect -2985 -957 -2973 -923
rect -3031 -972 -2973 -957
rect -2873 -787 -2815 -772
rect -2873 -821 -2861 -787
rect -2827 -821 -2815 -787
rect -2873 -855 -2815 -821
rect -2873 -889 -2861 -855
rect -2827 -889 -2815 -855
rect -2873 -923 -2815 -889
rect -2873 -957 -2861 -923
rect -2827 -957 -2815 -923
rect -2873 -972 -2815 -957
rect -2715 -787 -2657 -772
rect -2715 -821 -2703 -787
rect -2669 -821 -2657 -787
rect -2715 -855 -2657 -821
rect -2715 -889 -2703 -855
rect -2669 -889 -2657 -855
rect -2715 -923 -2657 -889
rect -2715 -957 -2703 -923
rect -2669 -957 -2657 -923
rect -2715 -972 -2657 -957
rect -2557 -787 -2499 -772
rect -2557 -821 -2545 -787
rect -2511 -821 -2499 -787
rect -2557 -855 -2499 -821
rect -2557 -889 -2545 -855
rect -2511 -889 -2499 -855
rect -2557 -923 -2499 -889
rect -2557 -957 -2545 -923
rect -2511 -957 -2499 -923
rect -2557 -972 -2499 -957
rect -2399 -787 -2341 -772
rect -2399 -821 -2387 -787
rect -2353 -821 -2341 -787
rect -2399 -855 -2341 -821
rect -2399 -889 -2387 -855
rect -2353 -889 -2341 -855
rect -2399 -923 -2341 -889
rect -2399 -957 -2387 -923
rect -2353 -957 -2341 -923
rect -2399 -972 -2341 -957
rect -2241 -787 -2183 -772
rect -2241 -821 -2229 -787
rect -2195 -821 -2183 -787
rect -2241 -855 -2183 -821
rect -2241 -889 -2229 -855
rect -2195 -889 -2183 -855
rect -2241 -923 -2183 -889
rect -2241 -957 -2229 -923
rect -2195 -957 -2183 -923
rect -2241 -972 -2183 -957
rect -2083 -787 -2025 -772
rect -2083 -821 -2071 -787
rect -2037 -821 -2025 -787
rect -2083 -855 -2025 -821
rect -2083 -889 -2071 -855
rect -2037 -889 -2025 -855
rect -2083 -923 -2025 -889
rect -2083 -957 -2071 -923
rect -2037 -957 -2025 -923
rect -2083 -972 -2025 -957
rect -1925 -787 -1867 -772
rect -1925 -821 -1913 -787
rect -1879 -821 -1867 -787
rect -1925 -855 -1867 -821
rect -1925 -889 -1913 -855
rect -1879 -889 -1867 -855
rect -1925 -923 -1867 -889
rect -1925 -957 -1913 -923
rect -1879 -957 -1867 -923
rect -1925 -972 -1867 -957
rect -1767 -787 -1709 -772
rect -1767 -821 -1755 -787
rect -1721 -821 -1709 -787
rect -1767 -855 -1709 -821
rect -1767 -889 -1755 -855
rect -1721 -889 -1709 -855
rect -1767 -923 -1709 -889
rect -1767 -957 -1755 -923
rect -1721 -957 -1709 -923
rect -1767 -972 -1709 -957
rect -1609 -787 -1551 -772
rect -1609 -821 -1597 -787
rect -1563 -821 -1551 -787
rect -1609 -855 -1551 -821
rect -1609 -889 -1597 -855
rect -1563 -889 -1551 -855
rect -1609 -923 -1551 -889
rect -1609 -957 -1597 -923
rect -1563 -957 -1551 -923
rect -1609 -972 -1551 -957
rect -1451 -787 -1393 -772
rect -1451 -821 -1439 -787
rect -1405 -821 -1393 -787
rect -1451 -855 -1393 -821
rect -1451 -889 -1439 -855
rect -1405 -889 -1393 -855
rect -1451 -923 -1393 -889
rect -1451 -957 -1439 -923
rect -1405 -957 -1393 -923
rect -1451 -972 -1393 -957
rect -1293 -787 -1235 -772
rect -1293 -821 -1281 -787
rect -1247 -821 -1235 -787
rect -1293 -855 -1235 -821
rect -1293 -889 -1281 -855
rect -1247 -889 -1235 -855
rect -1293 -923 -1235 -889
rect -1293 -957 -1281 -923
rect -1247 -957 -1235 -923
rect -1293 -972 -1235 -957
rect -1135 -787 -1077 -772
rect -1135 -821 -1123 -787
rect -1089 -821 -1077 -787
rect -1135 -855 -1077 -821
rect -1135 -889 -1123 -855
rect -1089 -889 -1077 -855
rect -1135 -923 -1077 -889
rect -1135 -957 -1123 -923
rect -1089 -957 -1077 -923
rect -1135 -972 -1077 -957
rect -977 -787 -919 -772
rect -977 -821 -965 -787
rect -931 -821 -919 -787
rect -977 -855 -919 -821
rect -977 -889 -965 -855
rect -931 -889 -919 -855
rect -977 -923 -919 -889
rect -977 -957 -965 -923
rect -931 -957 -919 -923
rect -977 -972 -919 -957
rect -819 -787 -761 -772
rect -819 -821 -807 -787
rect -773 -821 -761 -787
rect -819 -855 -761 -821
rect -819 -889 -807 -855
rect -773 -889 -761 -855
rect -819 -923 -761 -889
rect -819 -957 -807 -923
rect -773 -957 -761 -923
rect -819 -972 -761 -957
rect -661 -787 -603 -772
rect -661 -821 -649 -787
rect -615 -821 -603 -787
rect -661 -855 -603 -821
rect -661 -889 -649 -855
rect -615 -889 -603 -855
rect -661 -923 -603 -889
rect -661 -957 -649 -923
rect -615 -957 -603 -923
rect -661 -972 -603 -957
rect -503 -787 -445 -772
rect -503 -821 -491 -787
rect -457 -821 -445 -787
rect -503 -855 -445 -821
rect -503 -889 -491 -855
rect -457 -889 -445 -855
rect -503 -923 -445 -889
rect -503 -957 -491 -923
rect -457 -957 -445 -923
rect -503 -972 -445 -957
rect -345 -787 -287 -772
rect -345 -821 -333 -787
rect -299 -821 -287 -787
rect -345 -855 -287 -821
rect -345 -889 -333 -855
rect -299 -889 -287 -855
rect -345 -923 -287 -889
rect -345 -957 -333 -923
rect -299 -957 -287 -923
rect -345 -972 -287 -957
rect -187 -787 -129 -772
rect -187 -821 -175 -787
rect -141 -821 -129 -787
rect -187 -855 -129 -821
rect -187 -889 -175 -855
rect -141 -889 -129 -855
rect -187 -923 -129 -889
rect -187 -957 -175 -923
rect -141 -957 -129 -923
rect -187 -972 -129 -957
rect -29 -787 29 -772
rect -29 -821 -17 -787
rect 17 -821 29 -787
rect -29 -855 29 -821
rect -29 -889 -17 -855
rect 17 -889 29 -855
rect -29 -923 29 -889
rect -29 -957 -17 -923
rect 17 -957 29 -923
rect -29 -972 29 -957
rect 129 -787 187 -772
rect 129 -821 141 -787
rect 175 -821 187 -787
rect 129 -855 187 -821
rect 129 -889 141 -855
rect 175 -889 187 -855
rect 129 -923 187 -889
rect 129 -957 141 -923
rect 175 -957 187 -923
rect 129 -972 187 -957
rect 287 -787 345 -772
rect 287 -821 299 -787
rect 333 -821 345 -787
rect 287 -855 345 -821
rect 287 -889 299 -855
rect 333 -889 345 -855
rect 287 -923 345 -889
rect 287 -957 299 -923
rect 333 -957 345 -923
rect 287 -972 345 -957
rect 445 -787 503 -772
rect 445 -821 457 -787
rect 491 -821 503 -787
rect 445 -855 503 -821
rect 445 -889 457 -855
rect 491 -889 503 -855
rect 445 -923 503 -889
rect 445 -957 457 -923
rect 491 -957 503 -923
rect 445 -972 503 -957
rect 603 -787 661 -772
rect 603 -821 615 -787
rect 649 -821 661 -787
rect 603 -855 661 -821
rect 603 -889 615 -855
rect 649 -889 661 -855
rect 603 -923 661 -889
rect 603 -957 615 -923
rect 649 -957 661 -923
rect 603 -972 661 -957
rect 761 -787 819 -772
rect 761 -821 773 -787
rect 807 -821 819 -787
rect 761 -855 819 -821
rect 761 -889 773 -855
rect 807 -889 819 -855
rect 761 -923 819 -889
rect 761 -957 773 -923
rect 807 -957 819 -923
rect 761 -972 819 -957
rect 919 -787 977 -772
rect 919 -821 931 -787
rect 965 -821 977 -787
rect 919 -855 977 -821
rect 919 -889 931 -855
rect 965 -889 977 -855
rect 919 -923 977 -889
rect 919 -957 931 -923
rect 965 -957 977 -923
rect 919 -972 977 -957
rect 1077 -787 1135 -772
rect 1077 -821 1089 -787
rect 1123 -821 1135 -787
rect 1077 -855 1135 -821
rect 1077 -889 1089 -855
rect 1123 -889 1135 -855
rect 1077 -923 1135 -889
rect 1077 -957 1089 -923
rect 1123 -957 1135 -923
rect 1077 -972 1135 -957
rect 1235 -787 1293 -772
rect 1235 -821 1247 -787
rect 1281 -821 1293 -787
rect 1235 -855 1293 -821
rect 1235 -889 1247 -855
rect 1281 -889 1293 -855
rect 1235 -923 1293 -889
rect 1235 -957 1247 -923
rect 1281 -957 1293 -923
rect 1235 -972 1293 -957
rect 1393 -787 1451 -772
rect 1393 -821 1405 -787
rect 1439 -821 1451 -787
rect 1393 -855 1451 -821
rect 1393 -889 1405 -855
rect 1439 -889 1451 -855
rect 1393 -923 1451 -889
rect 1393 -957 1405 -923
rect 1439 -957 1451 -923
rect 1393 -972 1451 -957
rect 1551 -787 1609 -772
rect 1551 -821 1563 -787
rect 1597 -821 1609 -787
rect 1551 -855 1609 -821
rect 1551 -889 1563 -855
rect 1597 -889 1609 -855
rect 1551 -923 1609 -889
rect 1551 -957 1563 -923
rect 1597 -957 1609 -923
rect 1551 -972 1609 -957
rect 1709 -787 1767 -772
rect 1709 -821 1721 -787
rect 1755 -821 1767 -787
rect 1709 -855 1767 -821
rect 1709 -889 1721 -855
rect 1755 -889 1767 -855
rect 1709 -923 1767 -889
rect 1709 -957 1721 -923
rect 1755 -957 1767 -923
rect 1709 -972 1767 -957
rect 1867 -787 1925 -772
rect 1867 -821 1879 -787
rect 1913 -821 1925 -787
rect 1867 -855 1925 -821
rect 1867 -889 1879 -855
rect 1913 -889 1925 -855
rect 1867 -923 1925 -889
rect 1867 -957 1879 -923
rect 1913 -957 1925 -923
rect 1867 -972 1925 -957
rect 2025 -787 2083 -772
rect 2025 -821 2037 -787
rect 2071 -821 2083 -787
rect 2025 -855 2083 -821
rect 2025 -889 2037 -855
rect 2071 -889 2083 -855
rect 2025 -923 2083 -889
rect 2025 -957 2037 -923
rect 2071 -957 2083 -923
rect 2025 -972 2083 -957
rect 2183 -787 2241 -772
rect 2183 -821 2195 -787
rect 2229 -821 2241 -787
rect 2183 -855 2241 -821
rect 2183 -889 2195 -855
rect 2229 -889 2241 -855
rect 2183 -923 2241 -889
rect 2183 -957 2195 -923
rect 2229 -957 2241 -923
rect 2183 -972 2241 -957
rect 2341 -787 2399 -772
rect 2341 -821 2353 -787
rect 2387 -821 2399 -787
rect 2341 -855 2399 -821
rect 2341 -889 2353 -855
rect 2387 -889 2399 -855
rect 2341 -923 2399 -889
rect 2341 -957 2353 -923
rect 2387 -957 2399 -923
rect 2341 -972 2399 -957
rect 2499 -787 2557 -772
rect 2499 -821 2511 -787
rect 2545 -821 2557 -787
rect 2499 -855 2557 -821
rect 2499 -889 2511 -855
rect 2545 -889 2557 -855
rect 2499 -923 2557 -889
rect 2499 -957 2511 -923
rect 2545 -957 2557 -923
rect 2499 -972 2557 -957
rect 2657 -787 2715 -772
rect 2657 -821 2669 -787
rect 2703 -821 2715 -787
rect 2657 -855 2715 -821
rect 2657 -889 2669 -855
rect 2703 -889 2715 -855
rect 2657 -923 2715 -889
rect 2657 -957 2669 -923
rect 2703 -957 2715 -923
rect 2657 -972 2715 -957
rect 2815 -787 2873 -772
rect 2815 -821 2827 -787
rect 2861 -821 2873 -787
rect 2815 -855 2873 -821
rect 2815 -889 2827 -855
rect 2861 -889 2873 -855
rect 2815 -923 2873 -889
rect 2815 -957 2827 -923
rect 2861 -957 2873 -923
rect 2815 -972 2873 -957
rect 2973 -787 3031 -772
rect 2973 -821 2985 -787
rect 3019 -821 3031 -787
rect 2973 -855 3031 -821
rect 2973 -889 2985 -855
rect 3019 -889 3031 -855
rect 2973 -923 3031 -889
rect 2973 -957 2985 -923
rect 3019 -957 3031 -923
rect 2973 -972 3031 -957
rect 3131 -787 3189 -772
rect 3131 -821 3143 -787
rect 3177 -821 3189 -787
rect 3131 -855 3189 -821
rect 3131 -889 3143 -855
rect 3177 -889 3189 -855
rect 3131 -923 3189 -889
rect 3131 -957 3143 -923
rect 3177 -957 3189 -923
rect 3131 -972 3189 -957
<< mvpdiffc >>
rect -3177 923 -3143 957
rect -3177 855 -3143 889
rect -3177 787 -3143 821
rect -3019 923 -2985 957
rect -3019 855 -2985 889
rect -3019 787 -2985 821
rect -2861 923 -2827 957
rect -2861 855 -2827 889
rect -2861 787 -2827 821
rect -2703 923 -2669 957
rect -2703 855 -2669 889
rect -2703 787 -2669 821
rect -2545 923 -2511 957
rect -2545 855 -2511 889
rect -2545 787 -2511 821
rect -2387 923 -2353 957
rect -2387 855 -2353 889
rect -2387 787 -2353 821
rect -2229 923 -2195 957
rect -2229 855 -2195 889
rect -2229 787 -2195 821
rect -2071 923 -2037 957
rect -2071 855 -2037 889
rect -2071 787 -2037 821
rect -1913 923 -1879 957
rect -1913 855 -1879 889
rect -1913 787 -1879 821
rect -1755 923 -1721 957
rect -1755 855 -1721 889
rect -1755 787 -1721 821
rect -1597 923 -1563 957
rect -1597 855 -1563 889
rect -1597 787 -1563 821
rect -1439 923 -1405 957
rect -1439 855 -1405 889
rect -1439 787 -1405 821
rect -1281 923 -1247 957
rect -1281 855 -1247 889
rect -1281 787 -1247 821
rect -1123 923 -1089 957
rect -1123 855 -1089 889
rect -1123 787 -1089 821
rect -965 923 -931 957
rect -965 855 -931 889
rect -965 787 -931 821
rect -807 923 -773 957
rect -807 855 -773 889
rect -807 787 -773 821
rect -649 923 -615 957
rect -649 855 -615 889
rect -649 787 -615 821
rect -491 923 -457 957
rect -491 855 -457 889
rect -491 787 -457 821
rect -333 923 -299 957
rect -333 855 -299 889
rect -333 787 -299 821
rect -175 923 -141 957
rect -175 855 -141 889
rect -175 787 -141 821
rect -17 923 17 957
rect -17 855 17 889
rect -17 787 17 821
rect 141 923 175 957
rect 141 855 175 889
rect 141 787 175 821
rect 299 923 333 957
rect 299 855 333 889
rect 299 787 333 821
rect 457 923 491 957
rect 457 855 491 889
rect 457 787 491 821
rect 615 923 649 957
rect 615 855 649 889
rect 615 787 649 821
rect 773 923 807 957
rect 773 855 807 889
rect 773 787 807 821
rect 931 923 965 957
rect 931 855 965 889
rect 931 787 965 821
rect 1089 923 1123 957
rect 1089 855 1123 889
rect 1089 787 1123 821
rect 1247 923 1281 957
rect 1247 855 1281 889
rect 1247 787 1281 821
rect 1405 923 1439 957
rect 1405 855 1439 889
rect 1405 787 1439 821
rect 1563 923 1597 957
rect 1563 855 1597 889
rect 1563 787 1597 821
rect 1721 923 1755 957
rect 1721 855 1755 889
rect 1721 787 1755 821
rect 1879 923 1913 957
rect 1879 855 1913 889
rect 1879 787 1913 821
rect 2037 923 2071 957
rect 2037 855 2071 889
rect 2037 787 2071 821
rect 2195 923 2229 957
rect 2195 855 2229 889
rect 2195 787 2229 821
rect 2353 923 2387 957
rect 2353 855 2387 889
rect 2353 787 2387 821
rect 2511 923 2545 957
rect 2511 855 2545 889
rect 2511 787 2545 821
rect 2669 923 2703 957
rect 2669 855 2703 889
rect 2669 787 2703 821
rect 2827 923 2861 957
rect 2827 855 2861 889
rect 2827 787 2861 821
rect 2985 923 3019 957
rect 2985 855 3019 889
rect 2985 787 3019 821
rect 3143 923 3177 957
rect 3143 855 3177 889
rect 3143 787 3177 821
rect -3177 487 -3143 521
rect -3177 419 -3143 453
rect -3177 351 -3143 385
rect -3019 487 -2985 521
rect -3019 419 -2985 453
rect -3019 351 -2985 385
rect -2861 487 -2827 521
rect -2861 419 -2827 453
rect -2861 351 -2827 385
rect -2703 487 -2669 521
rect -2703 419 -2669 453
rect -2703 351 -2669 385
rect -2545 487 -2511 521
rect -2545 419 -2511 453
rect -2545 351 -2511 385
rect -2387 487 -2353 521
rect -2387 419 -2353 453
rect -2387 351 -2353 385
rect -2229 487 -2195 521
rect -2229 419 -2195 453
rect -2229 351 -2195 385
rect -2071 487 -2037 521
rect -2071 419 -2037 453
rect -2071 351 -2037 385
rect -1913 487 -1879 521
rect -1913 419 -1879 453
rect -1913 351 -1879 385
rect -1755 487 -1721 521
rect -1755 419 -1721 453
rect -1755 351 -1721 385
rect -1597 487 -1563 521
rect -1597 419 -1563 453
rect -1597 351 -1563 385
rect -1439 487 -1405 521
rect -1439 419 -1405 453
rect -1439 351 -1405 385
rect -1281 487 -1247 521
rect -1281 419 -1247 453
rect -1281 351 -1247 385
rect -1123 487 -1089 521
rect -1123 419 -1089 453
rect -1123 351 -1089 385
rect -965 487 -931 521
rect -965 419 -931 453
rect -965 351 -931 385
rect -807 487 -773 521
rect -807 419 -773 453
rect -807 351 -773 385
rect -649 487 -615 521
rect -649 419 -615 453
rect -649 351 -615 385
rect -491 487 -457 521
rect -491 419 -457 453
rect -491 351 -457 385
rect -333 487 -299 521
rect -333 419 -299 453
rect -333 351 -299 385
rect -175 487 -141 521
rect -175 419 -141 453
rect -175 351 -141 385
rect -17 487 17 521
rect -17 419 17 453
rect -17 351 17 385
rect 141 487 175 521
rect 141 419 175 453
rect 141 351 175 385
rect 299 487 333 521
rect 299 419 333 453
rect 299 351 333 385
rect 457 487 491 521
rect 457 419 491 453
rect 457 351 491 385
rect 615 487 649 521
rect 615 419 649 453
rect 615 351 649 385
rect 773 487 807 521
rect 773 419 807 453
rect 773 351 807 385
rect 931 487 965 521
rect 931 419 965 453
rect 931 351 965 385
rect 1089 487 1123 521
rect 1089 419 1123 453
rect 1089 351 1123 385
rect 1247 487 1281 521
rect 1247 419 1281 453
rect 1247 351 1281 385
rect 1405 487 1439 521
rect 1405 419 1439 453
rect 1405 351 1439 385
rect 1563 487 1597 521
rect 1563 419 1597 453
rect 1563 351 1597 385
rect 1721 487 1755 521
rect 1721 419 1755 453
rect 1721 351 1755 385
rect 1879 487 1913 521
rect 1879 419 1913 453
rect 1879 351 1913 385
rect 2037 487 2071 521
rect 2037 419 2071 453
rect 2037 351 2071 385
rect 2195 487 2229 521
rect 2195 419 2229 453
rect 2195 351 2229 385
rect 2353 487 2387 521
rect 2353 419 2387 453
rect 2353 351 2387 385
rect 2511 487 2545 521
rect 2511 419 2545 453
rect 2511 351 2545 385
rect 2669 487 2703 521
rect 2669 419 2703 453
rect 2669 351 2703 385
rect 2827 487 2861 521
rect 2827 419 2861 453
rect 2827 351 2861 385
rect 2985 487 3019 521
rect 2985 419 3019 453
rect 2985 351 3019 385
rect 3143 487 3177 521
rect 3143 419 3177 453
rect 3143 351 3177 385
rect -3177 51 -3143 85
rect -3177 -17 -3143 17
rect -3177 -85 -3143 -51
rect -3019 51 -2985 85
rect -3019 -17 -2985 17
rect -3019 -85 -2985 -51
rect -2861 51 -2827 85
rect -2861 -17 -2827 17
rect -2861 -85 -2827 -51
rect -2703 51 -2669 85
rect -2703 -17 -2669 17
rect -2703 -85 -2669 -51
rect -2545 51 -2511 85
rect -2545 -17 -2511 17
rect -2545 -85 -2511 -51
rect -2387 51 -2353 85
rect -2387 -17 -2353 17
rect -2387 -85 -2353 -51
rect -2229 51 -2195 85
rect -2229 -17 -2195 17
rect -2229 -85 -2195 -51
rect -2071 51 -2037 85
rect -2071 -17 -2037 17
rect -2071 -85 -2037 -51
rect -1913 51 -1879 85
rect -1913 -17 -1879 17
rect -1913 -85 -1879 -51
rect -1755 51 -1721 85
rect -1755 -17 -1721 17
rect -1755 -85 -1721 -51
rect -1597 51 -1563 85
rect -1597 -17 -1563 17
rect -1597 -85 -1563 -51
rect -1439 51 -1405 85
rect -1439 -17 -1405 17
rect -1439 -85 -1405 -51
rect -1281 51 -1247 85
rect -1281 -17 -1247 17
rect -1281 -85 -1247 -51
rect -1123 51 -1089 85
rect -1123 -17 -1089 17
rect -1123 -85 -1089 -51
rect -965 51 -931 85
rect -965 -17 -931 17
rect -965 -85 -931 -51
rect -807 51 -773 85
rect -807 -17 -773 17
rect -807 -85 -773 -51
rect -649 51 -615 85
rect -649 -17 -615 17
rect -649 -85 -615 -51
rect -491 51 -457 85
rect -491 -17 -457 17
rect -491 -85 -457 -51
rect -333 51 -299 85
rect -333 -17 -299 17
rect -333 -85 -299 -51
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect 299 51 333 85
rect 299 -17 333 17
rect 299 -85 333 -51
rect 457 51 491 85
rect 457 -17 491 17
rect 457 -85 491 -51
rect 615 51 649 85
rect 615 -17 649 17
rect 615 -85 649 -51
rect 773 51 807 85
rect 773 -17 807 17
rect 773 -85 807 -51
rect 931 51 965 85
rect 931 -17 965 17
rect 931 -85 965 -51
rect 1089 51 1123 85
rect 1089 -17 1123 17
rect 1089 -85 1123 -51
rect 1247 51 1281 85
rect 1247 -17 1281 17
rect 1247 -85 1281 -51
rect 1405 51 1439 85
rect 1405 -17 1439 17
rect 1405 -85 1439 -51
rect 1563 51 1597 85
rect 1563 -17 1597 17
rect 1563 -85 1597 -51
rect 1721 51 1755 85
rect 1721 -17 1755 17
rect 1721 -85 1755 -51
rect 1879 51 1913 85
rect 1879 -17 1913 17
rect 1879 -85 1913 -51
rect 2037 51 2071 85
rect 2037 -17 2071 17
rect 2037 -85 2071 -51
rect 2195 51 2229 85
rect 2195 -17 2229 17
rect 2195 -85 2229 -51
rect 2353 51 2387 85
rect 2353 -17 2387 17
rect 2353 -85 2387 -51
rect 2511 51 2545 85
rect 2511 -17 2545 17
rect 2511 -85 2545 -51
rect 2669 51 2703 85
rect 2669 -17 2703 17
rect 2669 -85 2703 -51
rect 2827 51 2861 85
rect 2827 -17 2861 17
rect 2827 -85 2861 -51
rect 2985 51 3019 85
rect 2985 -17 3019 17
rect 2985 -85 3019 -51
rect 3143 51 3177 85
rect 3143 -17 3177 17
rect 3143 -85 3177 -51
rect -3177 -385 -3143 -351
rect -3177 -453 -3143 -419
rect -3177 -521 -3143 -487
rect -3019 -385 -2985 -351
rect -3019 -453 -2985 -419
rect -3019 -521 -2985 -487
rect -2861 -385 -2827 -351
rect -2861 -453 -2827 -419
rect -2861 -521 -2827 -487
rect -2703 -385 -2669 -351
rect -2703 -453 -2669 -419
rect -2703 -521 -2669 -487
rect -2545 -385 -2511 -351
rect -2545 -453 -2511 -419
rect -2545 -521 -2511 -487
rect -2387 -385 -2353 -351
rect -2387 -453 -2353 -419
rect -2387 -521 -2353 -487
rect -2229 -385 -2195 -351
rect -2229 -453 -2195 -419
rect -2229 -521 -2195 -487
rect -2071 -385 -2037 -351
rect -2071 -453 -2037 -419
rect -2071 -521 -2037 -487
rect -1913 -385 -1879 -351
rect -1913 -453 -1879 -419
rect -1913 -521 -1879 -487
rect -1755 -385 -1721 -351
rect -1755 -453 -1721 -419
rect -1755 -521 -1721 -487
rect -1597 -385 -1563 -351
rect -1597 -453 -1563 -419
rect -1597 -521 -1563 -487
rect -1439 -385 -1405 -351
rect -1439 -453 -1405 -419
rect -1439 -521 -1405 -487
rect -1281 -385 -1247 -351
rect -1281 -453 -1247 -419
rect -1281 -521 -1247 -487
rect -1123 -385 -1089 -351
rect -1123 -453 -1089 -419
rect -1123 -521 -1089 -487
rect -965 -385 -931 -351
rect -965 -453 -931 -419
rect -965 -521 -931 -487
rect -807 -385 -773 -351
rect -807 -453 -773 -419
rect -807 -521 -773 -487
rect -649 -385 -615 -351
rect -649 -453 -615 -419
rect -649 -521 -615 -487
rect -491 -385 -457 -351
rect -491 -453 -457 -419
rect -491 -521 -457 -487
rect -333 -385 -299 -351
rect -333 -453 -299 -419
rect -333 -521 -299 -487
rect -175 -385 -141 -351
rect -175 -453 -141 -419
rect -175 -521 -141 -487
rect -17 -385 17 -351
rect -17 -453 17 -419
rect -17 -521 17 -487
rect 141 -385 175 -351
rect 141 -453 175 -419
rect 141 -521 175 -487
rect 299 -385 333 -351
rect 299 -453 333 -419
rect 299 -521 333 -487
rect 457 -385 491 -351
rect 457 -453 491 -419
rect 457 -521 491 -487
rect 615 -385 649 -351
rect 615 -453 649 -419
rect 615 -521 649 -487
rect 773 -385 807 -351
rect 773 -453 807 -419
rect 773 -521 807 -487
rect 931 -385 965 -351
rect 931 -453 965 -419
rect 931 -521 965 -487
rect 1089 -385 1123 -351
rect 1089 -453 1123 -419
rect 1089 -521 1123 -487
rect 1247 -385 1281 -351
rect 1247 -453 1281 -419
rect 1247 -521 1281 -487
rect 1405 -385 1439 -351
rect 1405 -453 1439 -419
rect 1405 -521 1439 -487
rect 1563 -385 1597 -351
rect 1563 -453 1597 -419
rect 1563 -521 1597 -487
rect 1721 -385 1755 -351
rect 1721 -453 1755 -419
rect 1721 -521 1755 -487
rect 1879 -385 1913 -351
rect 1879 -453 1913 -419
rect 1879 -521 1913 -487
rect 2037 -385 2071 -351
rect 2037 -453 2071 -419
rect 2037 -521 2071 -487
rect 2195 -385 2229 -351
rect 2195 -453 2229 -419
rect 2195 -521 2229 -487
rect 2353 -385 2387 -351
rect 2353 -453 2387 -419
rect 2353 -521 2387 -487
rect 2511 -385 2545 -351
rect 2511 -453 2545 -419
rect 2511 -521 2545 -487
rect 2669 -385 2703 -351
rect 2669 -453 2703 -419
rect 2669 -521 2703 -487
rect 2827 -385 2861 -351
rect 2827 -453 2861 -419
rect 2827 -521 2861 -487
rect 2985 -385 3019 -351
rect 2985 -453 3019 -419
rect 2985 -521 3019 -487
rect 3143 -385 3177 -351
rect 3143 -453 3177 -419
rect 3143 -521 3177 -487
rect -3177 -821 -3143 -787
rect -3177 -889 -3143 -855
rect -3177 -957 -3143 -923
rect -3019 -821 -2985 -787
rect -3019 -889 -2985 -855
rect -3019 -957 -2985 -923
rect -2861 -821 -2827 -787
rect -2861 -889 -2827 -855
rect -2861 -957 -2827 -923
rect -2703 -821 -2669 -787
rect -2703 -889 -2669 -855
rect -2703 -957 -2669 -923
rect -2545 -821 -2511 -787
rect -2545 -889 -2511 -855
rect -2545 -957 -2511 -923
rect -2387 -821 -2353 -787
rect -2387 -889 -2353 -855
rect -2387 -957 -2353 -923
rect -2229 -821 -2195 -787
rect -2229 -889 -2195 -855
rect -2229 -957 -2195 -923
rect -2071 -821 -2037 -787
rect -2071 -889 -2037 -855
rect -2071 -957 -2037 -923
rect -1913 -821 -1879 -787
rect -1913 -889 -1879 -855
rect -1913 -957 -1879 -923
rect -1755 -821 -1721 -787
rect -1755 -889 -1721 -855
rect -1755 -957 -1721 -923
rect -1597 -821 -1563 -787
rect -1597 -889 -1563 -855
rect -1597 -957 -1563 -923
rect -1439 -821 -1405 -787
rect -1439 -889 -1405 -855
rect -1439 -957 -1405 -923
rect -1281 -821 -1247 -787
rect -1281 -889 -1247 -855
rect -1281 -957 -1247 -923
rect -1123 -821 -1089 -787
rect -1123 -889 -1089 -855
rect -1123 -957 -1089 -923
rect -965 -821 -931 -787
rect -965 -889 -931 -855
rect -965 -957 -931 -923
rect -807 -821 -773 -787
rect -807 -889 -773 -855
rect -807 -957 -773 -923
rect -649 -821 -615 -787
rect -649 -889 -615 -855
rect -649 -957 -615 -923
rect -491 -821 -457 -787
rect -491 -889 -457 -855
rect -491 -957 -457 -923
rect -333 -821 -299 -787
rect -333 -889 -299 -855
rect -333 -957 -299 -923
rect -175 -821 -141 -787
rect -175 -889 -141 -855
rect -175 -957 -141 -923
rect -17 -821 17 -787
rect -17 -889 17 -855
rect -17 -957 17 -923
rect 141 -821 175 -787
rect 141 -889 175 -855
rect 141 -957 175 -923
rect 299 -821 333 -787
rect 299 -889 333 -855
rect 299 -957 333 -923
rect 457 -821 491 -787
rect 457 -889 491 -855
rect 457 -957 491 -923
rect 615 -821 649 -787
rect 615 -889 649 -855
rect 615 -957 649 -923
rect 773 -821 807 -787
rect 773 -889 807 -855
rect 773 -957 807 -923
rect 931 -821 965 -787
rect 931 -889 965 -855
rect 931 -957 965 -923
rect 1089 -821 1123 -787
rect 1089 -889 1123 -855
rect 1089 -957 1123 -923
rect 1247 -821 1281 -787
rect 1247 -889 1281 -855
rect 1247 -957 1281 -923
rect 1405 -821 1439 -787
rect 1405 -889 1439 -855
rect 1405 -957 1439 -923
rect 1563 -821 1597 -787
rect 1563 -889 1597 -855
rect 1563 -957 1597 -923
rect 1721 -821 1755 -787
rect 1721 -889 1755 -855
rect 1721 -957 1755 -923
rect 1879 -821 1913 -787
rect 1879 -889 1913 -855
rect 1879 -957 1913 -923
rect 2037 -821 2071 -787
rect 2037 -889 2071 -855
rect 2037 -957 2071 -923
rect 2195 -821 2229 -787
rect 2195 -889 2229 -855
rect 2195 -957 2229 -923
rect 2353 -821 2387 -787
rect 2353 -889 2387 -855
rect 2353 -957 2387 -923
rect 2511 -821 2545 -787
rect 2511 -889 2545 -855
rect 2511 -957 2545 -923
rect 2669 -821 2703 -787
rect 2669 -889 2703 -855
rect 2669 -957 2703 -923
rect 2827 -821 2861 -787
rect 2827 -889 2861 -855
rect 2827 -957 2861 -923
rect 2985 -821 3019 -787
rect 2985 -889 3019 -855
rect 2985 -957 3019 -923
rect 3143 -821 3177 -787
rect 3143 -889 3177 -855
rect 3143 -957 3177 -923
<< mvnsubdiff >>
rect -3323 1191 3323 1203
rect -3323 1157 -3213 1191
rect -3179 1157 -3145 1191
rect -3111 1157 -3077 1191
rect -3043 1157 -3009 1191
rect -2975 1157 -2941 1191
rect -2907 1157 -2873 1191
rect -2839 1157 -2805 1191
rect -2771 1157 -2737 1191
rect -2703 1157 -2669 1191
rect -2635 1157 -2601 1191
rect -2567 1157 -2533 1191
rect -2499 1157 -2465 1191
rect -2431 1157 -2397 1191
rect -2363 1157 -2329 1191
rect -2295 1157 -2261 1191
rect -2227 1157 -2193 1191
rect -2159 1157 -2125 1191
rect -2091 1157 -2057 1191
rect -2023 1157 -1989 1191
rect -1955 1157 -1921 1191
rect -1887 1157 -1853 1191
rect -1819 1157 -1785 1191
rect -1751 1157 -1717 1191
rect -1683 1157 -1649 1191
rect -1615 1157 -1581 1191
rect -1547 1157 -1513 1191
rect -1479 1157 -1445 1191
rect -1411 1157 -1377 1191
rect -1343 1157 -1309 1191
rect -1275 1157 -1241 1191
rect -1207 1157 -1173 1191
rect -1139 1157 -1105 1191
rect -1071 1157 -1037 1191
rect -1003 1157 -969 1191
rect -935 1157 -901 1191
rect -867 1157 -833 1191
rect -799 1157 -765 1191
rect -731 1157 -697 1191
rect -663 1157 -629 1191
rect -595 1157 -561 1191
rect -527 1157 -493 1191
rect -459 1157 -425 1191
rect -391 1157 -357 1191
rect -323 1157 -289 1191
rect -255 1157 -221 1191
rect -187 1157 -153 1191
rect -119 1157 -85 1191
rect -51 1157 -17 1191
rect 17 1157 51 1191
rect 85 1157 119 1191
rect 153 1157 187 1191
rect 221 1157 255 1191
rect 289 1157 323 1191
rect 357 1157 391 1191
rect 425 1157 459 1191
rect 493 1157 527 1191
rect 561 1157 595 1191
rect 629 1157 663 1191
rect 697 1157 731 1191
rect 765 1157 799 1191
rect 833 1157 867 1191
rect 901 1157 935 1191
rect 969 1157 1003 1191
rect 1037 1157 1071 1191
rect 1105 1157 1139 1191
rect 1173 1157 1207 1191
rect 1241 1157 1275 1191
rect 1309 1157 1343 1191
rect 1377 1157 1411 1191
rect 1445 1157 1479 1191
rect 1513 1157 1547 1191
rect 1581 1157 1615 1191
rect 1649 1157 1683 1191
rect 1717 1157 1751 1191
rect 1785 1157 1819 1191
rect 1853 1157 1887 1191
rect 1921 1157 1955 1191
rect 1989 1157 2023 1191
rect 2057 1157 2091 1191
rect 2125 1157 2159 1191
rect 2193 1157 2227 1191
rect 2261 1157 2295 1191
rect 2329 1157 2363 1191
rect 2397 1157 2431 1191
rect 2465 1157 2499 1191
rect 2533 1157 2567 1191
rect 2601 1157 2635 1191
rect 2669 1157 2703 1191
rect 2737 1157 2771 1191
rect 2805 1157 2839 1191
rect 2873 1157 2907 1191
rect 2941 1157 2975 1191
rect 3009 1157 3043 1191
rect 3077 1157 3111 1191
rect 3145 1157 3179 1191
rect 3213 1157 3323 1191
rect -3323 1145 3323 1157
rect -3323 1071 -3265 1145
rect -3323 1037 -3311 1071
rect -3277 1037 -3265 1071
rect 3265 1071 3323 1145
rect -3323 1003 -3265 1037
rect -3323 969 -3311 1003
rect -3277 969 -3265 1003
rect 3265 1037 3277 1071
rect 3311 1037 3323 1071
rect 3265 1003 3323 1037
rect -3323 935 -3265 969
rect -3323 901 -3311 935
rect -3277 901 -3265 935
rect -3323 867 -3265 901
rect -3323 833 -3311 867
rect -3277 833 -3265 867
rect -3323 799 -3265 833
rect -3323 765 -3311 799
rect -3277 765 -3265 799
rect 3265 969 3277 1003
rect 3311 969 3323 1003
rect 3265 935 3323 969
rect 3265 901 3277 935
rect 3311 901 3323 935
rect 3265 867 3323 901
rect 3265 833 3277 867
rect 3311 833 3323 867
rect 3265 799 3323 833
rect -3323 731 -3265 765
rect -3323 697 -3311 731
rect -3277 697 -3265 731
rect -3323 663 -3265 697
rect 3265 765 3277 799
rect 3311 765 3323 799
rect 3265 731 3323 765
rect 3265 697 3277 731
rect 3311 697 3323 731
rect -3323 629 -3311 663
rect -3277 629 -3265 663
rect 3265 663 3323 697
rect -3323 595 -3265 629
rect -3323 561 -3311 595
rect -3277 561 -3265 595
rect -3323 527 -3265 561
rect 3265 629 3277 663
rect 3311 629 3323 663
rect 3265 595 3323 629
rect 3265 561 3277 595
rect 3311 561 3323 595
rect -3323 493 -3311 527
rect -3277 493 -3265 527
rect -3323 459 -3265 493
rect -3323 425 -3311 459
rect -3277 425 -3265 459
rect -3323 391 -3265 425
rect -3323 357 -3311 391
rect -3277 357 -3265 391
rect -3323 323 -3265 357
rect 3265 527 3323 561
rect 3265 493 3277 527
rect 3311 493 3323 527
rect 3265 459 3323 493
rect 3265 425 3277 459
rect 3311 425 3323 459
rect 3265 391 3323 425
rect 3265 357 3277 391
rect 3311 357 3323 391
rect -3323 289 -3311 323
rect -3277 289 -3265 323
rect -3323 255 -3265 289
rect -3323 221 -3311 255
rect -3277 221 -3265 255
rect 3265 323 3323 357
rect 3265 289 3277 323
rect 3311 289 3323 323
rect 3265 255 3323 289
rect -3323 187 -3265 221
rect 3265 221 3277 255
rect 3311 221 3323 255
rect -3323 153 -3311 187
rect -3277 153 -3265 187
rect -3323 119 -3265 153
rect -3323 85 -3311 119
rect -3277 85 -3265 119
rect 3265 187 3323 221
rect 3265 153 3277 187
rect 3311 153 3323 187
rect 3265 119 3323 153
rect -3323 51 -3265 85
rect -3323 17 -3311 51
rect -3277 17 -3265 51
rect -3323 -17 -3265 17
rect -3323 -51 -3311 -17
rect -3277 -51 -3265 -17
rect -3323 -85 -3265 -51
rect -3323 -119 -3311 -85
rect -3277 -119 -3265 -85
rect 3265 85 3277 119
rect 3311 85 3323 119
rect 3265 51 3323 85
rect 3265 17 3277 51
rect 3311 17 3323 51
rect 3265 -17 3323 17
rect 3265 -51 3277 -17
rect 3311 -51 3323 -17
rect 3265 -85 3323 -51
rect -3323 -153 -3265 -119
rect -3323 -187 -3311 -153
rect -3277 -187 -3265 -153
rect -3323 -221 -3265 -187
rect 3265 -119 3277 -85
rect 3311 -119 3323 -85
rect 3265 -153 3323 -119
rect 3265 -187 3277 -153
rect 3311 -187 3323 -153
rect -3323 -255 -3311 -221
rect -3277 -255 -3265 -221
rect 3265 -221 3323 -187
rect -3323 -289 -3265 -255
rect -3323 -323 -3311 -289
rect -3277 -323 -3265 -289
rect -3323 -357 -3265 -323
rect 3265 -255 3277 -221
rect 3311 -255 3323 -221
rect 3265 -289 3323 -255
rect 3265 -323 3277 -289
rect 3311 -323 3323 -289
rect -3323 -391 -3311 -357
rect -3277 -391 -3265 -357
rect -3323 -425 -3265 -391
rect -3323 -459 -3311 -425
rect -3277 -459 -3265 -425
rect -3323 -493 -3265 -459
rect -3323 -527 -3311 -493
rect -3277 -527 -3265 -493
rect -3323 -561 -3265 -527
rect 3265 -357 3323 -323
rect 3265 -391 3277 -357
rect 3311 -391 3323 -357
rect 3265 -425 3323 -391
rect 3265 -459 3277 -425
rect 3311 -459 3323 -425
rect 3265 -493 3323 -459
rect 3265 -527 3277 -493
rect 3311 -527 3323 -493
rect -3323 -595 -3311 -561
rect -3277 -595 -3265 -561
rect -3323 -629 -3265 -595
rect -3323 -663 -3311 -629
rect -3277 -663 -3265 -629
rect 3265 -561 3323 -527
rect 3265 -595 3277 -561
rect 3311 -595 3323 -561
rect 3265 -629 3323 -595
rect -3323 -697 -3265 -663
rect 3265 -663 3277 -629
rect 3311 -663 3323 -629
rect -3323 -731 -3311 -697
rect -3277 -731 -3265 -697
rect -3323 -765 -3265 -731
rect -3323 -799 -3311 -765
rect -3277 -799 -3265 -765
rect 3265 -697 3323 -663
rect 3265 -731 3277 -697
rect 3311 -731 3323 -697
rect 3265 -765 3323 -731
rect -3323 -833 -3265 -799
rect -3323 -867 -3311 -833
rect -3277 -867 -3265 -833
rect -3323 -901 -3265 -867
rect -3323 -935 -3311 -901
rect -3277 -935 -3265 -901
rect -3323 -969 -3265 -935
rect -3323 -1003 -3311 -969
rect -3277 -1003 -3265 -969
rect 3265 -799 3277 -765
rect 3311 -799 3323 -765
rect 3265 -833 3323 -799
rect 3265 -867 3277 -833
rect 3311 -867 3323 -833
rect 3265 -901 3323 -867
rect 3265 -935 3277 -901
rect 3311 -935 3323 -901
rect 3265 -969 3323 -935
rect -3323 -1037 -3265 -1003
rect -3323 -1071 -3311 -1037
rect -3277 -1071 -3265 -1037
rect 3265 -1003 3277 -969
rect 3311 -1003 3323 -969
rect 3265 -1037 3323 -1003
rect -3323 -1145 -3265 -1071
rect 3265 -1071 3277 -1037
rect 3311 -1071 3323 -1037
rect 3265 -1145 3323 -1071
rect -3323 -1157 3323 -1145
rect -3323 -1191 -3213 -1157
rect -3179 -1191 -3145 -1157
rect -3111 -1191 -3077 -1157
rect -3043 -1191 -3009 -1157
rect -2975 -1191 -2941 -1157
rect -2907 -1191 -2873 -1157
rect -2839 -1191 -2805 -1157
rect -2771 -1191 -2737 -1157
rect -2703 -1191 -2669 -1157
rect -2635 -1191 -2601 -1157
rect -2567 -1191 -2533 -1157
rect -2499 -1191 -2465 -1157
rect -2431 -1191 -2397 -1157
rect -2363 -1191 -2329 -1157
rect -2295 -1191 -2261 -1157
rect -2227 -1191 -2193 -1157
rect -2159 -1191 -2125 -1157
rect -2091 -1191 -2057 -1157
rect -2023 -1191 -1989 -1157
rect -1955 -1191 -1921 -1157
rect -1887 -1191 -1853 -1157
rect -1819 -1191 -1785 -1157
rect -1751 -1191 -1717 -1157
rect -1683 -1191 -1649 -1157
rect -1615 -1191 -1581 -1157
rect -1547 -1191 -1513 -1157
rect -1479 -1191 -1445 -1157
rect -1411 -1191 -1377 -1157
rect -1343 -1191 -1309 -1157
rect -1275 -1191 -1241 -1157
rect -1207 -1191 -1173 -1157
rect -1139 -1191 -1105 -1157
rect -1071 -1191 -1037 -1157
rect -1003 -1191 -969 -1157
rect -935 -1191 -901 -1157
rect -867 -1191 -833 -1157
rect -799 -1191 -765 -1157
rect -731 -1191 -697 -1157
rect -663 -1191 -629 -1157
rect -595 -1191 -561 -1157
rect -527 -1191 -493 -1157
rect -459 -1191 -425 -1157
rect -391 -1191 -357 -1157
rect -323 -1191 -289 -1157
rect -255 -1191 -221 -1157
rect -187 -1191 -153 -1157
rect -119 -1191 -85 -1157
rect -51 -1191 -17 -1157
rect 17 -1191 51 -1157
rect 85 -1191 119 -1157
rect 153 -1191 187 -1157
rect 221 -1191 255 -1157
rect 289 -1191 323 -1157
rect 357 -1191 391 -1157
rect 425 -1191 459 -1157
rect 493 -1191 527 -1157
rect 561 -1191 595 -1157
rect 629 -1191 663 -1157
rect 697 -1191 731 -1157
rect 765 -1191 799 -1157
rect 833 -1191 867 -1157
rect 901 -1191 935 -1157
rect 969 -1191 1003 -1157
rect 1037 -1191 1071 -1157
rect 1105 -1191 1139 -1157
rect 1173 -1191 1207 -1157
rect 1241 -1191 1275 -1157
rect 1309 -1191 1343 -1157
rect 1377 -1191 1411 -1157
rect 1445 -1191 1479 -1157
rect 1513 -1191 1547 -1157
rect 1581 -1191 1615 -1157
rect 1649 -1191 1683 -1157
rect 1717 -1191 1751 -1157
rect 1785 -1191 1819 -1157
rect 1853 -1191 1887 -1157
rect 1921 -1191 1955 -1157
rect 1989 -1191 2023 -1157
rect 2057 -1191 2091 -1157
rect 2125 -1191 2159 -1157
rect 2193 -1191 2227 -1157
rect 2261 -1191 2295 -1157
rect 2329 -1191 2363 -1157
rect 2397 -1191 2431 -1157
rect 2465 -1191 2499 -1157
rect 2533 -1191 2567 -1157
rect 2601 -1191 2635 -1157
rect 2669 -1191 2703 -1157
rect 2737 -1191 2771 -1157
rect 2805 -1191 2839 -1157
rect 2873 -1191 2907 -1157
rect 2941 -1191 2975 -1157
rect 3009 -1191 3043 -1157
rect 3077 -1191 3111 -1157
rect 3145 -1191 3179 -1157
rect 3213 -1191 3323 -1157
rect -3323 -1203 3323 -1191
<< mvnsubdiffcont >>
rect -3213 1157 -3179 1191
rect -3145 1157 -3111 1191
rect -3077 1157 -3043 1191
rect -3009 1157 -2975 1191
rect -2941 1157 -2907 1191
rect -2873 1157 -2839 1191
rect -2805 1157 -2771 1191
rect -2737 1157 -2703 1191
rect -2669 1157 -2635 1191
rect -2601 1157 -2567 1191
rect -2533 1157 -2499 1191
rect -2465 1157 -2431 1191
rect -2397 1157 -2363 1191
rect -2329 1157 -2295 1191
rect -2261 1157 -2227 1191
rect -2193 1157 -2159 1191
rect -2125 1157 -2091 1191
rect -2057 1157 -2023 1191
rect -1989 1157 -1955 1191
rect -1921 1157 -1887 1191
rect -1853 1157 -1819 1191
rect -1785 1157 -1751 1191
rect -1717 1157 -1683 1191
rect -1649 1157 -1615 1191
rect -1581 1157 -1547 1191
rect -1513 1157 -1479 1191
rect -1445 1157 -1411 1191
rect -1377 1157 -1343 1191
rect -1309 1157 -1275 1191
rect -1241 1157 -1207 1191
rect -1173 1157 -1139 1191
rect -1105 1157 -1071 1191
rect -1037 1157 -1003 1191
rect -969 1157 -935 1191
rect -901 1157 -867 1191
rect -833 1157 -799 1191
rect -765 1157 -731 1191
rect -697 1157 -663 1191
rect -629 1157 -595 1191
rect -561 1157 -527 1191
rect -493 1157 -459 1191
rect -425 1157 -391 1191
rect -357 1157 -323 1191
rect -289 1157 -255 1191
rect -221 1157 -187 1191
rect -153 1157 -119 1191
rect -85 1157 -51 1191
rect -17 1157 17 1191
rect 51 1157 85 1191
rect 119 1157 153 1191
rect 187 1157 221 1191
rect 255 1157 289 1191
rect 323 1157 357 1191
rect 391 1157 425 1191
rect 459 1157 493 1191
rect 527 1157 561 1191
rect 595 1157 629 1191
rect 663 1157 697 1191
rect 731 1157 765 1191
rect 799 1157 833 1191
rect 867 1157 901 1191
rect 935 1157 969 1191
rect 1003 1157 1037 1191
rect 1071 1157 1105 1191
rect 1139 1157 1173 1191
rect 1207 1157 1241 1191
rect 1275 1157 1309 1191
rect 1343 1157 1377 1191
rect 1411 1157 1445 1191
rect 1479 1157 1513 1191
rect 1547 1157 1581 1191
rect 1615 1157 1649 1191
rect 1683 1157 1717 1191
rect 1751 1157 1785 1191
rect 1819 1157 1853 1191
rect 1887 1157 1921 1191
rect 1955 1157 1989 1191
rect 2023 1157 2057 1191
rect 2091 1157 2125 1191
rect 2159 1157 2193 1191
rect 2227 1157 2261 1191
rect 2295 1157 2329 1191
rect 2363 1157 2397 1191
rect 2431 1157 2465 1191
rect 2499 1157 2533 1191
rect 2567 1157 2601 1191
rect 2635 1157 2669 1191
rect 2703 1157 2737 1191
rect 2771 1157 2805 1191
rect 2839 1157 2873 1191
rect 2907 1157 2941 1191
rect 2975 1157 3009 1191
rect 3043 1157 3077 1191
rect 3111 1157 3145 1191
rect 3179 1157 3213 1191
rect -3311 1037 -3277 1071
rect -3311 969 -3277 1003
rect 3277 1037 3311 1071
rect -3311 901 -3277 935
rect -3311 833 -3277 867
rect -3311 765 -3277 799
rect 3277 969 3311 1003
rect 3277 901 3311 935
rect 3277 833 3311 867
rect -3311 697 -3277 731
rect 3277 765 3311 799
rect 3277 697 3311 731
rect -3311 629 -3277 663
rect -3311 561 -3277 595
rect 3277 629 3311 663
rect 3277 561 3311 595
rect -3311 493 -3277 527
rect -3311 425 -3277 459
rect -3311 357 -3277 391
rect 3277 493 3311 527
rect 3277 425 3311 459
rect 3277 357 3311 391
rect -3311 289 -3277 323
rect -3311 221 -3277 255
rect 3277 289 3311 323
rect 3277 221 3311 255
rect -3311 153 -3277 187
rect -3311 85 -3277 119
rect 3277 153 3311 187
rect -3311 17 -3277 51
rect -3311 -51 -3277 -17
rect -3311 -119 -3277 -85
rect 3277 85 3311 119
rect 3277 17 3311 51
rect 3277 -51 3311 -17
rect -3311 -187 -3277 -153
rect 3277 -119 3311 -85
rect 3277 -187 3311 -153
rect -3311 -255 -3277 -221
rect -3311 -323 -3277 -289
rect 3277 -255 3311 -221
rect 3277 -323 3311 -289
rect -3311 -391 -3277 -357
rect -3311 -459 -3277 -425
rect -3311 -527 -3277 -493
rect 3277 -391 3311 -357
rect 3277 -459 3311 -425
rect 3277 -527 3311 -493
rect -3311 -595 -3277 -561
rect -3311 -663 -3277 -629
rect 3277 -595 3311 -561
rect 3277 -663 3311 -629
rect -3311 -731 -3277 -697
rect -3311 -799 -3277 -765
rect 3277 -731 3311 -697
rect -3311 -867 -3277 -833
rect -3311 -935 -3277 -901
rect -3311 -1003 -3277 -969
rect 3277 -799 3311 -765
rect 3277 -867 3311 -833
rect 3277 -935 3311 -901
rect -3311 -1071 -3277 -1037
rect 3277 -1003 3311 -969
rect 3277 -1071 3311 -1037
rect -3213 -1191 -3179 -1157
rect -3145 -1191 -3111 -1157
rect -3077 -1191 -3043 -1157
rect -3009 -1191 -2975 -1157
rect -2941 -1191 -2907 -1157
rect -2873 -1191 -2839 -1157
rect -2805 -1191 -2771 -1157
rect -2737 -1191 -2703 -1157
rect -2669 -1191 -2635 -1157
rect -2601 -1191 -2567 -1157
rect -2533 -1191 -2499 -1157
rect -2465 -1191 -2431 -1157
rect -2397 -1191 -2363 -1157
rect -2329 -1191 -2295 -1157
rect -2261 -1191 -2227 -1157
rect -2193 -1191 -2159 -1157
rect -2125 -1191 -2091 -1157
rect -2057 -1191 -2023 -1157
rect -1989 -1191 -1955 -1157
rect -1921 -1191 -1887 -1157
rect -1853 -1191 -1819 -1157
rect -1785 -1191 -1751 -1157
rect -1717 -1191 -1683 -1157
rect -1649 -1191 -1615 -1157
rect -1581 -1191 -1547 -1157
rect -1513 -1191 -1479 -1157
rect -1445 -1191 -1411 -1157
rect -1377 -1191 -1343 -1157
rect -1309 -1191 -1275 -1157
rect -1241 -1191 -1207 -1157
rect -1173 -1191 -1139 -1157
rect -1105 -1191 -1071 -1157
rect -1037 -1191 -1003 -1157
rect -969 -1191 -935 -1157
rect -901 -1191 -867 -1157
rect -833 -1191 -799 -1157
rect -765 -1191 -731 -1157
rect -697 -1191 -663 -1157
rect -629 -1191 -595 -1157
rect -561 -1191 -527 -1157
rect -493 -1191 -459 -1157
rect -425 -1191 -391 -1157
rect -357 -1191 -323 -1157
rect -289 -1191 -255 -1157
rect -221 -1191 -187 -1157
rect -153 -1191 -119 -1157
rect -85 -1191 -51 -1157
rect -17 -1191 17 -1157
rect 51 -1191 85 -1157
rect 119 -1191 153 -1157
rect 187 -1191 221 -1157
rect 255 -1191 289 -1157
rect 323 -1191 357 -1157
rect 391 -1191 425 -1157
rect 459 -1191 493 -1157
rect 527 -1191 561 -1157
rect 595 -1191 629 -1157
rect 663 -1191 697 -1157
rect 731 -1191 765 -1157
rect 799 -1191 833 -1157
rect 867 -1191 901 -1157
rect 935 -1191 969 -1157
rect 1003 -1191 1037 -1157
rect 1071 -1191 1105 -1157
rect 1139 -1191 1173 -1157
rect 1207 -1191 1241 -1157
rect 1275 -1191 1309 -1157
rect 1343 -1191 1377 -1157
rect 1411 -1191 1445 -1157
rect 1479 -1191 1513 -1157
rect 1547 -1191 1581 -1157
rect 1615 -1191 1649 -1157
rect 1683 -1191 1717 -1157
rect 1751 -1191 1785 -1157
rect 1819 -1191 1853 -1157
rect 1887 -1191 1921 -1157
rect 1955 -1191 1989 -1157
rect 2023 -1191 2057 -1157
rect 2091 -1191 2125 -1157
rect 2159 -1191 2193 -1157
rect 2227 -1191 2261 -1157
rect 2295 -1191 2329 -1157
rect 2363 -1191 2397 -1157
rect 2431 -1191 2465 -1157
rect 2499 -1191 2533 -1157
rect 2567 -1191 2601 -1157
rect 2635 -1191 2669 -1157
rect 2703 -1191 2737 -1157
rect 2771 -1191 2805 -1157
rect 2839 -1191 2873 -1157
rect 2907 -1191 2941 -1157
rect 2975 -1191 3009 -1157
rect 3043 -1191 3077 -1157
rect 3111 -1191 3145 -1157
rect 3179 -1191 3213 -1157
<< poly >>
rect -3131 1053 -3031 1069
rect -3131 1019 -3098 1053
rect -3064 1019 -3031 1053
rect -3131 972 -3031 1019
rect -2973 1053 -2873 1069
rect -2973 1019 -2940 1053
rect -2906 1019 -2873 1053
rect -2973 972 -2873 1019
rect -2815 1053 -2715 1069
rect -2815 1019 -2782 1053
rect -2748 1019 -2715 1053
rect -2815 972 -2715 1019
rect -2657 1053 -2557 1069
rect -2657 1019 -2624 1053
rect -2590 1019 -2557 1053
rect -2657 972 -2557 1019
rect -2499 1053 -2399 1069
rect -2499 1019 -2466 1053
rect -2432 1019 -2399 1053
rect -2499 972 -2399 1019
rect -2341 1053 -2241 1069
rect -2341 1019 -2308 1053
rect -2274 1019 -2241 1053
rect -2341 972 -2241 1019
rect -2183 1053 -2083 1069
rect -2183 1019 -2150 1053
rect -2116 1019 -2083 1053
rect -2183 972 -2083 1019
rect -2025 1053 -1925 1069
rect -2025 1019 -1992 1053
rect -1958 1019 -1925 1053
rect -2025 972 -1925 1019
rect -1867 1053 -1767 1069
rect -1867 1019 -1834 1053
rect -1800 1019 -1767 1053
rect -1867 972 -1767 1019
rect -1709 1053 -1609 1069
rect -1709 1019 -1676 1053
rect -1642 1019 -1609 1053
rect -1709 972 -1609 1019
rect -1551 1053 -1451 1069
rect -1551 1019 -1518 1053
rect -1484 1019 -1451 1053
rect -1551 972 -1451 1019
rect -1393 1053 -1293 1069
rect -1393 1019 -1360 1053
rect -1326 1019 -1293 1053
rect -1393 972 -1293 1019
rect -1235 1053 -1135 1069
rect -1235 1019 -1202 1053
rect -1168 1019 -1135 1053
rect -1235 972 -1135 1019
rect -1077 1053 -977 1069
rect -1077 1019 -1044 1053
rect -1010 1019 -977 1053
rect -1077 972 -977 1019
rect -919 1053 -819 1069
rect -919 1019 -886 1053
rect -852 1019 -819 1053
rect -919 972 -819 1019
rect -761 1053 -661 1069
rect -761 1019 -728 1053
rect -694 1019 -661 1053
rect -761 972 -661 1019
rect -603 1053 -503 1069
rect -603 1019 -570 1053
rect -536 1019 -503 1053
rect -603 972 -503 1019
rect -445 1053 -345 1069
rect -445 1019 -412 1053
rect -378 1019 -345 1053
rect -445 972 -345 1019
rect -287 1053 -187 1069
rect -287 1019 -254 1053
rect -220 1019 -187 1053
rect -287 972 -187 1019
rect -129 1053 -29 1069
rect -129 1019 -96 1053
rect -62 1019 -29 1053
rect -129 972 -29 1019
rect 29 1053 129 1069
rect 29 1019 62 1053
rect 96 1019 129 1053
rect 29 972 129 1019
rect 187 1053 287 1069
rect 187 1019 220 1053
rect 254 1019 287 1053
rect 187 972 287 1019
rect 345 1053 445 1069
rect 345 1019 378 1053
rect 412 1019 445 1053
rect 345 972 445 1019
rect 503 1053 603 1069
rect 503 1019 536 1053
rect 570 1019 603 1053
rect 503 972 603 1019
rect 661 1053 761 1069
rect 661 1019 694 1053
rect 728 1019 761 1053
rect 661 972 761 1019
rect 819 1053 919 1069
rect 819 1019 852 1053
rect 886 1019 919 1053
rect 819 972 919 1019
rect 977 1053 1077 1069
rect 977 1019 1010 1053
rect 1044 1019 1077 1053
rect 977 972 1077 1019
rect 1135 1053 1235 1069
rect 1135 1019 1168 1053
rect 1202 1019 1235 1053
rect 1135 972 1235 1019
rect 1293 1053 1393 1069
rect 1293 1019 1326 1053
rect 1360 1019 1393 1053
rect 1293 972 1393 1019
rect 1451 1053 1551 1069
rect 1451 1019 1484 1053
rect 1518 1019 1551 1053
rect 1451 972 1551 1019
rect 1609 1053 1709 1069
rect 1609 1019 1642 1053
rect 1676 1019 1709 1053
rect 1609 972 1709 1019
rect 1767 1053 1867 1069
rect 1767 1019 1800 1053
rect 1834 1019 1867 1053
rect 1767 972 1867 1019
rect 1925 1053 2025 1069
rect 1925 1019 1958 1053
rect 1992 1019 2025 1053
rect 1925 972 2025 1019
rect 2083 1053 2183 1069
rect 2083 1019 2116 1053
rect 2150 1019 2183 1053
rect 2083 972 2183 1019
rect 2241 1053 2341 1069
rect 2241 1019 2274 1053
rect 2308 1019 2341 1053
rect 2241 972 2341 1019
rect 2399 1053 2499 1069
rect 2399 1019 2432 1053
rect 2466 1019 2499 1053
rect 2399 972 2499 1019
rect 2557 1053 2657 1069
rect 2557 1019 2590 1053
rect 2624 1019 2657 1053
rect 2557 972 2657 1019
rect 2715 1053 2815 1069
rect 2715 1019 2748 1053
rect 2782 1019 2815 1053
rect 2715 972 2815 1019
rect 2873 1053 2973 1069
rect 2873 1019 2906 1053
rect 2940 1019 2973 1053
rect 2873 972 2973 1019
rect 3031 1053 3131 1069
rect 3031 1019 3064 1053
rect 3098 1019 3131 1053
rect 3031 972 3131 1019
rect -3131 725 -3031 772
rect -3131 691 -3098 725
rect -3064 691 -3031 725
rect -3131 675 -3031 691
rect -2973 725 -2873 772
rect -2973 691 -2940 725
rect -2906 691 -2873 725
rect -2973 675 -2873 691
rect -2815 725 -2715 772
rect -2815 691 -2782 725
rect -2748 691 -2715 725
rect -2815 675 -2715 691
rect -2657 725 -2557 772
rect -2657 691 -2624 725
rect -2590 691 -2557 725
rect -2657 675 -2557 691
rect -2499 725 -2399 772
rect -2499 691 -2466 725
rect -2432 691 -2399 725
rect -2499 675 -2399 691
rect -2341 725 -2241 772
rect -2341 691 -2308 725
rect -2274 691 -2241 725
rect -2341 675 -2241 691
rect -2183 725 -2083 772
rect -2183 691 -2150 725
rect -2116 691 -2083 725
rect -2183 675 -2083 691
rect -2025 725 -1925 772
rect -2025 691 -1992 725
rect -1958 691 -1925 725
rect -2025 675 -1925 691
rect -1867 725 -1767 772
rect -1867 691 -1834 725
rect -1800 691 -1767 725
rect -1867 675 -1767 691
rect -1709 725 -1609 772
rect -1709 691 -1676 725
rect -1642 691 -1609 725
rect -1709 675 -1609 691
rect -1551 725 -1451 772
rect -1551 691 -1518 725
rect -1484 691 -1451 725
rect -1551 675 -1451 691
rect -1393 725 -1293 772
rect -1393 691 -1360 725
rect -1326 691 -1293 725
rect -1393 675 -1293 691
rect -1235 725 -1135 772
rect -1235 691 -1202 725
rect -1168 691 -1135 725
rect -1235 675 -1135 691
rect -1077 725 -977 772
rect -1077 691 -1044 725
rect -1010 691 -977 725
rect -1077 675 -977 691
rect -919 725 -819 772
rect -919 691 -886 725
rect -852 691 -819 725
rect -919 675 -819 691
rect -761 725 -661 772
rect -761 691 -728 725
rect -694 691 -661 725
rect -761 675 -661 691
rect -603 725 -503 772
rect -603 691 -570 725
rect -536 691 -503 725
rect -603 675 -503 691
rect -445 725 -345 772
rect -445 691 -412 725
rect -378 691 -345 725
rect -445 675 -345 691
rect -287 725 -187 772
rect -287 691 -254 725
rect -220 691 -187 725
rect -287 675 -187 691
rect -129 725 -29 772
rect -129 691 -96 725
rect -62 691 -29 725
rect -129 675 -29 691
rect 29 725 129 772
rect 29 691 62 725
rect 96 691 129 725
rect 29 675 129 691
rect 187 725 287 772
rect 187 691 220 725
rect 254 691 287 725
rect 187 675 287 691
rect 345 725 445 772
rect 345 691 378 725
rect 412 691 445 725
rect 345 675 445 691
rect 503 725 603 772
rect 503 691 536 725
rect 570 691 603 725
rect 503 675 603 691
rect 661 725 761 772
rect 661 691 694 725
rect 728 691 761 725
rect 661 675 761 691
rect 819 725 919 772
rect 819 691 852 725
rect 886 691 919 725
rect 819 675 919 691
rect 977 725 1077 772
rect 977 691 1010 725
rect 1044 691 1077 725
rect 977 675 1077 691
rect 1135 725 1235 772
rect 1135 691 1168 725
rect 1202 691 1235 725
rect 1135 675 1235 691
rect 1293 725 1393 772
rect 1293 691 1326 725
rect 1360 691 1393 725
rect 1293 675 1393 691
rect 1451 725 1551 772
rect 1451 691 1484 725
rect 1518 691 1551 725
rect 1451 675 1551 691
rect 1609 725 1709 772
rect 1609 691 1642 725
rect 1676 691 1709 725
rect 1609 675 1709 691
rect 1767 725 1867 772
rect 1767 691 1800 725
rect 1834 691 1867 725
rect 1767 675 1867 691
rect 1925 725 2025 772
rect 1925 691 1958 725
rect 1992 691 2025 725
rect 1925 675 2025 691
rect 2083 725 2183 772
rect 2083 691 2116 725
rect 2150 691 2183 725
rect 2083 675 2183 691
rect 2241 725 2341 772
rect 2241 691 2274 725
rect 2308 691 2341 725
rect 2241 675 2341 691
rect 2399 725 2499 772
rect 2399 691 2432 725
rect 2466 691 2499 725
rect 2399 675 2499 691
rect 2557 725 2657 772
rect 2557 691 2590 725
rect 2624 691 2657 725
rect 2557 675 2657 691
rect 2715 725 2815 772
rect 2715 691 2748 725
rect 2782 691 2815 725
rect 2715 675 2815 691
rect 2873 725 2973 772
rect 2873 691 2906 725
rect 2940 691 2973 725
rect 2873 675 2973 691
rect 3031 725 3131 772
rect 3031 691 3064 725
rect 3098 691 3131 725
rect 3031 675 3131 691
rect -3131 617 -3031 633
rect -3131 583 -3098 617
rect -3064 583 -3031 617
rect -3131 536 -3031 583
rect -2973 617 -2873 633
rect -2973 583 -2940 617
rect -2906 583 -2873 617
rect -2973 536 -2873 583
rect -2815 617 -2715 633
rect -2815 583 -2782 617
rect -2748 583 -2715 617
rect -2815 536 -2715 583
rect -2657 617 -2557 633
rect -2657 583 -2624 617
rect -2590 583 -2557 617
rect -2657 536 -2557 583
rect -2499 617 -2399 633
rect -2499 583 -2466 617
rect -2432 583 -2399 617
rect -2499 536 -2399 583
rect -2341 617 -2241 633
rect -2341 583 -2308 617
rect -2274 583 -2241 617
rect -2341 536 -2241 583
rect -2183 617 -2083 633
rect -2183 583 -2150 617
rect -2116 583 -2083 617
rect -2183 536 -2083 583
rect -2025 617 -1925 633
rect -2025 583 -1992 617
rect -1958 583 -1925 617
rect -2025 536 -1925 583
rect -1867 617 -1767 633
rect -1867 583 -1834 617
rect -1800 583 -1767 617
rect -1867 536 -1767 583
rect -1709 617 -1609 633
rect -1709 583 -1676 617
rect -1642 583 -1609 617
rect -1709 536 -1609 583
rect -1551 617 -1451 633
rect -1551 583 -1518 617
rect -1484 583 -1451 617
rect -1551 536 -1451 583
rect -1393 617 -1293 633
rect -1393 583 -1360 617
rect -1326 583 -1293 617
rect -1393 536 -1293 583
rect -1235 617 -1135 633
rect -1235 583 -1202 617
rect -1168 583 -1135 617
rect -1235 536 -1135 583
rect -1077 617 -977 633
rect -1077 583 -1044 617
rect -1010 583 -977 617
rect -1077 536 -977 583
rect -919 617 -819 633
rect -919 583 -886 617
rect -852 583 -819 617
rect -919 536 -819 583
rect -761 617 -661 633
rect -761 583 -728 617
rect -694 583 -661 617
rect -761 536 -661 583
rect -603 617 -503 633
rect -603 583 -570 617
rect -536 583 -503 617
rect -603 536 -503 583
rect -445 617 -345 633
rect -445 583 -412 617
rect -378 583 -345 617
rect -445 536 -345 583
rect -287 617 -187 633
rect -287 583 -254 617
rect -220 583 -187 617
rect -287 536 -187 583
rect -129 617 -29 633
rect -129 583 -96 617
rect -62 583 -29 617
rect -129 536 -29 583
rect 29 617 129 633
rect 29 583 62 617
rect 96 583 129 617
rect 29 536 129 583
rect 187 617 287 633
rect 187 583 220 617
rect 254 583 287 617
rect 187 536 287 583
rect 345 617 445 633
rect 345 583 378 617
rect 412 583 445 617
rect 345 536 445 583
rect 503 617 603 633
rect 503 583 536 617
rect 570 583 603 617
rect 503 536 603 583
rect 661 617 761 633
rect 661 583 694 617
rect 728 583 761 617
rect 661 536 761 583
rect 819 617 919 633
rect 819 583 852 617
rect 886 583 919 617
rect 819 536 919 583
rect 977 617 1077 633
rect 977 583 1010 617
rect 1044 583 1077 617
rect 977 536 1077 583
rect 1135 617 1235 633
rect 1135 583 1168 617
rect 1202 583 1235 617
rect 1135 536 1235 583
rect 1293 617 1393 633
rect 1293 583 1326 617
rect 1360 583 1393 617
rect 1293 536 1393 583
rect 1451 617 1551 633
rect 1451 583 1484 617
rect 1518 583 1551 617
rect 1451 536 1551 583
rect 1609 617 1709 633
rect 1609 583 1642 617
rect 1676 583 1709 617
rect 1609 536 1709 583
rect 1767 617 1867 633
rect 1767 583 1800 617
rect 1834 583 1867 617
rect 1767 536 1867 583
rect 1925 617 2025 633
rect 1925 583 1958 617
rect 1992 583 2025 617
rect 1925 536 2025 583
rect 2083 617 2183 633
rect 2083 583 2116 617
rect 2150 583 2183 617
rect 2083 536 2183 583
rect 2241 617 2341 633
rect 2241 583 2274 617
rect 2308 583 2341 617
rect 2241 536 2341 583
rect 2399 617 2499 633
rect 2399 583 2432 617
rect 2466 583 2499 617
rect 2399 536 2499 583
rect 2557 617 2657 633
rect 2557 583 2590 617
rect 2624 583 2657 617
rect 2557 536 2657 583
rect 2715 617 2815 633
rect 2715 583 2748 617
rect 2782 583 2815 617
rect 2715 536 2815 583
rect 2873 617 2973 633
rect 2873 583 2906 617
rect 2940 583 2973 617
rect 2873 536 2973 583
rect 3031 617 3131 633
rect 3031 583 3064 617
rect 3098 583 3131 617
rect 3031 536 3131 583
rect -3131 289 -3031 336
rect -3131 255 -3098 289
rect -3064 255 -3031 289
rect -3131 239 -3031 255
rect -2973 289 -2873 336
rect -2973 255 -2940 289
rect -2906 255 -2873 289
rect -2973 239 -2873 255
rect -2815 289 -2715 336
rect -2815 255 -2782 289
rect -2748 255 -2715 289
rect -2815 239 -2715 255
rect -2657 289 -2557 336
rect -2657 255 -2624 289
rect -2590 255 -2557 289
rect -2657 239 -2557 255
rect -2499 289 -2399 336
rect -2499 255 -2466 289
rect -2432 255 -2399 289
rect -2499 239 -2399 255
rect -2341 289 -2241 336
rect -2341 255 -2308 289
rect -2274 255 -2241 289
rect -2341 239 -2241 255
rect -2183 289 -2083 336
rect -2183 255 -2150 289
rect -2116 255 -2083 289
rect -2183 239 -2083 255
rect -2025 289 -1925 336
rect -2025 255 -1992 289
rect -1958 255 -1925 289
rect -2025 239 -1925 255
rect -1867 289 -1767 336
rect -1867 255 -1834 289
rect -1800 255 -1767 289
rect -1867 239 -1767 255
rect -1709 289 -1609 336
rect -1709 255 -1676 289
rect -1642 255 -1609 289
rect -1709 239 -1609 255
rect -1551 289 -1451 336
rect -1551 255 -1518 289
rect -1484 255 -1451 289
rect -1551 239 -1451 255
rect -1393 289 -1293 336
rect -1393 255 -1360 289
rect -1326 255 -1293 289
rect -1393 239 -1293 255
rect -1235 289 -1135 336
rect -1235 255 -1202 289
rect -1168 255 -1135 289
rect -1235 239 -1135 255
rect -1077 289 -977 336
rect -1077 255 -1044 289
rect -1010 255 -977 289
rect -1077 239 -977 255
rect -919 289 -819 336
rect -919 255 -886 289
rect -852 255 -819 289
rect -919 239 -819 255
rect -761 289 -661 336
rect -761 255 -728 289
rect -694 255 -661 289
rect -761 239 -661 255
rect -603 289 -503 336
rect -603 255 -570 289
rect -536 255 -503 289
rect -603 239 -503 255
rect -445 289 -345 336
rect -445 255 -412 289
rect -378 255 -345 289
rect -445 239 -345 255
rect -287 289 -187 336
rect -287 255 -254 289
rect -220 255 -187 289
rect -287 239 -187 255
rect -129 289 -29 336
rect -129 255 -96 289
rect -62 255 -29 289
rect -129 239 -29 255
rect 29 289 129 336
rect 29 255 62 289
rect 96 255 129 289
rect 29 239 129 255
rect 187 289 287 336
rect 187 255 220 289
rect 254 255 287 289
rect 187 239 287 255
rect 345 289 445 336
rect 345 255 378 289
rect 412 255 445 289
rect 345 239 445 255
rect 503 289 603 336
rect 503 255 536 289
rect 570 255 603 289
rect 503 239 603 255
rect 661 289 761 336
rect 661 255 694 289
rect 728 255 761 289
rect 661 239 761 255
rect 819 289 919 336
rect 819 255 852 289
rect 886 255 919 289
rect 819 239 919 255
rect 977 289 1077 336
rect 977 255 1010 289
rect 1044 255 1077 289
rect 977 239 1077 255
rect 1135 289 1235 336
rect 1135 255 1168 289
rect 1202 255 1235 289
rect 1135 239 1235 255
rect 1293 289 1393 336
rect 1293 255 1326 289
rect 1360 255 1393 289
rect 1293 239 1393 255
rect 1451 289 1551 336
rect 1451 255 1484 289
rect 1518 255 1551 289
rect 1451 239 1551 255
rect 1609 289 1709 336
rect 1609 255 1642 289
rect 1676 255 1709 289
rect 1609 239 1709 255
rect 1767 289 1867 336
rect 1767 255 1800 289
rect 1834 255 1867 289
rect 1767 239 1867 255
rect 1925 289 2025 336
rect 1925 255 1958 289
rect 1992 255 2025 289
rect 1925 239 2025 255
rect 2083 289 2183 336
rect 2083 255 2116 289
rect 2150 255 2183 289
rect 2083 239 2183 255
rect 2241 289 2341 336
rect 2241 255 2274 289
rect 2308 255 2341 289
rect 2241 239 2341 255
rect 2399 289 2499 336
rect 2399 255 2432 289
rect 2466 255 2499 289
rect 2399 239 2499 255
rect 2557 289 2657 336
rect 2557 255 2590 289
rect 2624 255 2657 289
rect 2557 239 2657 255
rect 2715 289 2815 336
rect 2715 255 2748 289
rect 2782 255 2815 289
rect 2715 239 2815 255
rect 2873 289 2973 336
rect 2873 255 2906 289
rect 2940 255 2973 289
rect 2873 239 2973 255
rect 3031 289 3131 336
rect 3031 255 3064 289
rect 3098 255 3131 289
rect 3031 239 3131 255
rect -3131 181 -3031 197
rect -3131 147 -3098 181
rect -3064 147 -3031 181
rect -3131 100 -3031 147
rect -2973 181 -2873 197
rect -2973 147 -2940 181
rect -2906 147 -2873 181
rect -2973 100 -2873 147
rect -2815 181 -2715 197
rect -2815 147 -2782 181
rect -2748 147 -2715 181
rect -2815 100 -2715 147
rect -2657 181 -2557 197
rect -2657 147 -2624 181
rect -2590 147 -2557 181
rect -2657 100 -2557 147
rect -2499 181 -2399 197
rect -2499 147 -2466 181
rect -2432 147 -2399 181
rect -2499 100 -2399 147
rect -2341 181 -2241 197
rect -2341 147 -2308 181
rect -2274 147 -2241 181
rect -2341 100 -2241 147
rect -2183 181 -2083 197
rect -2183 147 -2150 181
rect -2116 147 -2083 181
rect -2183 100 -2083 147
rect -2025 181 -1925 197
rect -2025 147 -1992 181
rect -1958 147 -1925 181
rect -2025 100 -1925 147
rect -1867 181 -1767 197
rect -1867 147 -1834 181
rect -1800 147 -1767 181
rect -1867 100 -1767 147
rect -1709 181 -1609 197
rect -1709 147 -1676 181
rect -1642 147 -1609 181
rect -1709 100 -1609 147
rect -1551 181 -1451 197
rect -1551 147 -1518 181
rect -1484 147 -1451 181
rect -1551 100 -1451 147
rect -1393 181 -1293 197
rect -1393 147 -1360 181
rect -1326 147 -1293 181
rect -1393 100 -1293 147
rect -1235 181 -1135 197
rect -1235 147 -1202 181
rect -1168 147 -1135 181
rect -1235 100 -1135 147
rect -1077 181 -977 197
rect -1077 147 -1044 181
rect -1010 147 -977 181
rect -1077 100 -977 147
rect -919 181 -819 197
rect -919 147 -886 181
rect -852 147 -819 181
rect -919 100 -819 147
rect -761 181 -661 197
rect -761 147 -728 181
rect -694 147 -661 181
rect -761 100 -661 147
rect -603 181 -503 197
rect -603 147 -570 181
rect -536 147 -503 181
rect -603 100 -503 147
rect -445 181 -345 197
rect -445 147 -412 181
rect -378 147 -345 181
rect -445 100 -345 147
rect -287 181 -187 197
rect -287 147 -254 181
rect -220 147 -187 181
rect -287 100 -187 147
rect -129 181 -29 197
rect -129 147 -96 181
rect -62 147 -29 181
rect -129 100 -29 147
rect 29 181 129 197
rect 29 147 62 181
rect 96 147 129 181
rect 29 100 129 147
rect 187 181 287 197
rect 187 147 220 181
rect 254 147 287 181
rect 187 100 287 147
rect 345 181 445 197
rect 345 147 378 181
rect 412 147 445 181
rect 345 100 445 147
rect 503 181 603 197
rect 503 147 536 181
rect 570 147 603 181
rect 503 100 603 147
rect 661 181 761 197
rect 661 147 694 181
rect 728 147 761 181
rect 661 100 761 147
rect 819 181 919 197
rect 819 147 852 181
rect 886 147 919 181
rect 819 100 919 147
rect 977 181 1077 197
rect 977 147 1010 181
rect 1044 147 1077 181
rect 977 100 1077 147
rect 1135 181 1235 197
rect 1135 147 1168 181
rect 1202 147 1235 181
rect 1135 100 1235 147
rect 1293 181 1393 197
rect 1293 147 1326 181
rect 1360 147 1393 181
rect 1293 100 1393 147
rect 1451 181 1551 197
rect 1451 147 1484 181
rect 1518 147 1551 181
rect 1451 100 1551 147
rect 1609 181 1709 197
rect 1609 147 1642 181
rect 1676 147 1709 181
rect 1609 100 1709 147
rect 1767 181 1867 197
rect 1767 147 1800 181
rect 1834 147 1867 181
rect 1767 100 1867 147
rect 1925 181 2025 197
rect 1925 147 1958 181
rect 1992 147 2025 181
rect 1925 100 2025 147
rect 2083 181 2183 197
rect 2083 147 2116 181
rect 2150 147 2183 181
rect 2083 100 2183 147
rect 2241 181 2341 197
rect 2241 147 2274 181
rect 2308 147 2341 181
rect 2241 100 2341 147
rect 2399 181 2499 197
rect 2399 147 2432 181
rect 2466 147 2499 181
rect 2399 100 2499 147
rect 2557 181 2657 197
rect 2557 147 2590 181
rect 2624 147 2657 181
rect 2557 100 2657 147
rect 2715 181 2815 197
rect 2715 147 2748 181
rect 2782 147 2815 181
rect 2715 100 2815 147
rect 2873 181 2973 197
rect 2873 147 2906 181
rect 2940 147 2973 181
rect 2873 100 2973 147
rect 3031 181 3131 197
rect 3031 147 3064 181
rect 3098 147 3131 181
rect 3031 100 3131 147
rect -3131 -147 -3031 -100
rect -3131 -181 -3098 -147
rect -3064 -181 -3031 -147
rect -3131 -197 -3031 -181
rect -2973 -147 -2873 -100
rect -2973 -181 -2940 -147
rect -2906 -181 -2873 -147
rect -2973 -197 -2873 -181
rect -2815 -147 -2715 -100
rect -2815 -181 -2782 -147
rect -2748 -181 -2715 -147
rect -2815 -197 -2715 -181
rect -2657 -147 -2557 -100
rect -2657 -181 -2624 -147
rect -2590 -181 -2557 -147
rect -2657 -197 -2557 -181
rect -2499 -147 -2399 -100
rect -2499 -181 -2466 -147
rect -2432 -181 -2399 -147
rect -2499 -197 -2399 -181
rect -2341 -147 -2241 -100
rect -2341 -181 -2308 -147
rect -2274 -181 -2241 -147
rect -2341 -197 -2241 -181
rect -2183 -147 -2083 -100
rect -2183 -181 -2150 -147
rect -2116 -181 -2083 -147
rect -2183 -197 -2083 -181
rect -2025 -147 -1925 -100
rect -2025 -181 -1992 -147
rect -1958 -181 -1925 -147
rect -2025 -197 -1925 -181
rect -1867 -147 -1767 -100
rect -1867 -181 -1834 -147
rect -1800 -181 -1767 -147
rect -1867 -197 -1767 -181
rect -1709 -147 -1609 -100
rect -1709 -181 -1676 -147
rect -1642 -181 -1609 -147
rect -1709 -197 -1609 -181
rect -1551 -147 -1451 -100
rect -1551 -181 -1518 -147
rect -1484 -181 -1451 -147
rect -1551 -197 -1451 -181
rect -1393 -147 -1293 -100
rect -1393 -181 -1360 -147
rect -1326 -181 -1293 -147
rect -1393 -197 -1293 -181
rect -1235 -147 -1135 -100
rect -1235 -181 -1202 -147
rect -1168 -181 -1135 -147
rect -1235 -197 -1135 -181
rect -1077 -147 -977 -100
rect -1077 -181 -1044 -147
rect -1010 -181 -977 -147
rect -1077 -197 -977 -181
rect -919 -147 -819 -100
rect -919 -181 -886 -147
rect -852 -181 -819 -147
rect -919 -197 -819 -181
rect -761 -147 -661 -100
rect -761 -181 -728 -147
rect -694 -181 -661 -147
rect -761 -197 -661 -181
rect -603 -147 -503 -100
rect -603 -181 -570 -147
rect -536 -181 -503 -147
rect -603 -197 -503 -181
rect -445 -147 -345 -100
rect -445 -181 -412 -147
rect -378 -181 -345 -147
rect -445 -197 -345 -181
rect -287 -147 -187 -100
rect -287 -181 -254 -147
rect -220 -181 -187 -147
rect -287 -197 -187 -181
rect -129 -147 -29 -100
rect -129 -181 -96 -147
rect -62 -181 -29 -147
rect -129 -197 -29 -181
rect 29 -147 129 -100
rect 29 -181 62 -147
rect 96 -181 129 -147
rect 29 -197 129 -181
rect 187 -147 287 -100
rect 187 -181 220 -147
rect 254 -181 287 -147
rect 187 -197 287 -181
rect 345 -147 445 -100
rect 345 -181 378 -147
rect 412 -181 445 -147
rect 345 -197 445 -181
rect 503 -147 603 -100
rect 503 -181 536 -147
rect 570 -181 603 -147
rect 503 -197 603 -181
rect 661 -147 761 -100
rect 661 -181 694 -147
rect 728 -181 761 -147
rect 661 -197 761 -181
rect 819 -147 919 -100
rect 819 -181 852 -147
rect 886 -181 919 -147
rect 819 -197 919 -181
rect 977 -147 1077 -100
rect 977 -181 1010 -147
rect 1044 -181 1077 -147
rect 977 -197 1077 -181
rect 1135 -147 1235 -100
rect 1135 -181 1168 -147
rect 1202 -181 1235 -147
rect 1135 -197 1235 -181
rect 1293 -147 1393 -100
rect 1293 -181 1326 -147
rect 1360 -181 1393 -147
rect 1293 -197 1393 -181
rect 1451 -147 1551 -100
rect 1451 -181 1484 -147
rect 1518 -181 1551 -147
rect 1451 -197 1551 -181
rect 1609 -147 1709 -100
rect 1609 -181 1642 -147
rect 1676 -181 1709 -147
rect 1609 -197 1709 -181
rect 1767 -147 1867 -100
rect 1767 -181 1800 -147
rect 1834 -181 1867 -147
rect 1767 -197 1867 -181
rect 1925 -147 2025 -100
rect 1925 -181 1958 -147
rect 1992 -181 2025 -147
rect 1925 -197 2025 -181
rect 2083 -147 2183 -100
rect 2083 -181 2116 -147
rect 2150 -181 2183 -147
rect 2083 -197 2183 -181
rect 2241 -147 2341 -100
rect 2241 -181 2274 -147
rect 2308 -181 2341 -147
rect 2241 -197 2341 -181
rect 2399 -147 2499 -100
rect 2399 -181 2432 -147
rect 2466 -181 2499 -147
rect 2399 -197 2499 -181
rect 2557 -147 2657 -100
rect 2557 -181 2590 -147
rect 2624 -181 2657 -147
rect 2557 -197 2657 -181
rect 2715 -147 2815 -100
rect 2715 -181 2748 -147
rect 2782 -181 2815 -147
rect 2715 -197 2815 -181
rect 2873 -147 2973 -100
rect 2873 -181 2906 -147
rect 2940 -181 2973 -147
rect 2873 -197 2973 -181
rect 3031 -147 3131 -100
rect 3031 -181 3064 -147
rect 3098 -181 3131 -147
rect 3031 -197 3131 -181
rect -3131 -255 -3031 -239
rect -3131 -289 -3098 -255
rect -3064 -289 -3031 -255
rect -3131 -336 -3031 -289
rect -2973 -255 -2873 -239
rect -2973 -289 -2940 -255
rect -2906 -289 -2873 -255
rect -2973 -336 -2873 -289
rect -2815 -255 -2715 -239
rect -2815 -289 -2782 -255
rect -2748 -289 -2715 -255
rect -2815 -336 -2715 -289
rect -2657 -255 -2557 -239
rect -2657 -289 -2624 -255
rect -2590 -289 -2557 -255
rect -2657 -336 -2557 -289
rect -2499 -255 -2399 -239
rect -2499 -289 -2466 -255
rect -2432 -289 -2399 -255
rect -2499 -336 -2399 -289
rect -2341 -255 -2241 -239
rect -2341 -289 -2308 -255
rect -2274 -289 -2241 -255
rect -2341 -336 -2241 -289
rect -2183 -255 -2083 -239
rect -2183 -289 -2150 -255
rect -2116 -289 -2083 -255
rect -2183 -336 -2083 -289
rect -2025 -255 -1925 -239
rect -2025 -289 -1992 -255
rect -1958 -289 -1925 -255
rect -2025 -336 -1925 -289
rect -1867 -255 -1767 -239
rect -1867 -289 -1834 -255
rect -1800 -289 -1767 -255
rect -1867 -336 -1767 -289
rect -1709 -255 -1609 -239
rect -1709 -289 -1676 -255
rect -1642 -289 -1609 -255
rect -1709 -336 -1609 -289
rect -1551 -255 -1451 -239
rect -1551 -289 -1518 -255
rect -1484 -289 -1451 -255
rect -1551 -336 -1451 -289
rect -1393 -255 -1293 -239
rect -1393 -289 -1360 -255
rect -1326 -289 -1293 -255
rect -1393 -336 -1293 -289
rect -1235 -255 -1135 -239
rect -1235 -289 -1202 -255
rect -1168 -289 -1135 -255
rect -1235 -336 -1135 -289
rect -1077 -255 -977 -239
rect -1077 -289 -1044 -255
rect -1010 -289 -977 -255
rect -1077 -336 -977 -289
rect -919 -255 -819 -239
rect -919 -289 -886 -255
rect -852 -289 -819 -255
rect -919 -336 -819 -289
rect -761 -255 -661 -239
rect -761 -289 -728 -255
rect -694 -289 -661 -255
rect -761 -336 -661 -289
rect -603 -255 -503 -239
rect -603 -289 -570 -255
rect -536 -289 -503 -255
rect -603 -336 -503 -289
rect -445 -255 -345 -239
rect -445 -289 -412 -255
rect -378 -289 -345 -255
rect -445 -336 -345 -289
rect -287 -255 -187 -239
rect -287 -289 -254 -255
rect -220 -289 -187 -255
rect -287 -336 -187 -289
rect -129 -255 -29 -239
rect -129 -289 -96 -255
rect -62 -289 -29 -255
rect -129 -336 -29 -289
rect 29 -255 129 -239
rect 29 -289 62 -255
rect 96 -289 129 -255
rect 29 -336 129 -289
rect 187 -255 287 -239
rect 187 -289 220 -255
rect 254 -289 287 -255
rect 187 -336 287 -289
rect 345 -255 445 -239
rect 345 -289 378 -255
rect 412 -289 445 -255
rect 345 -336 445 -289
rect 503 -255 603 -239
rect 503 -289 536 -255
rect 570 -289 603 -255
rect 503 -336 603 -289
rect 661 -255 761 -239
rect 661 -289 694 -255
rect 728 -289 761 -255
rect 661 -336 761 -289
rect 819 -255 919 -239
rect 819 -289 852 -255
rect 886 -289 919 -255
rect 819 -336 919 -289
rect 977 -255 1077 -239
rect 977 -289 1010 -255
rect 1044 -289 1077 -255
rect 977 -336 1077 -289
rect 1135 -255 1235 -239
rect 1135 -289 1168 -255
rect 1202 -289 1235 -255
rect 1135 -336 1235 -289
rect 1293 -255 1393 -239
rect 1293 -289 1326 -255
rect 1360 -289 1393 -255
rect 1293 -336 1393 -289
rect 1451 -255 1551 -239
rect 1451 -289 1484 -255
rect 1518 -289 1551 -255
rect 1451 -336 1551 -289
rect 1609 -255 1709 -239
rect 1609 -289 1642 -255
rect 1676 -289 1709 -255
rect 1609 -336 1709 -289
rect 1767 -255 1867 -239
rect 1767 -289 1800 -255
rect 1834 -289 1867 -255
rect 1767 -336 1867 -289
rect 1925 -255 2025 -239
rect 1925 -289 1958 -255
rect 1992 -289 2025 -255
rect 1925 -336 2025 -289
rect 2083 -255 2183 -239
rect 2083 -289 2116 -255
rect 2150 -289 2183 -255
rect 2083 -336 2183 -289
rect 2241 -255 2341 -239
rect 2241 -289 2274 -255
rect 2308 -289 2341 -255
rect 2241 -336 2341 -289
rect 2399 -255 2499 -239
rect 2399 -289 2432 -255
rect 2466 -289 2499 -255
rect 2399 -336 2499 -289
rect 2557 -255 2657 -239
rect 2557 -289 2590 -255
rect 2624 -289 2657 -255
rect 2557 -336 2657 -289
rect 2715 -255 2815 -239
rect 2715 -289 2748 -255
rect 2782 -289 2815 -255
rect 2715 -336 2815 -289
rect 2873 -255 2973 -239
rect 2873 -289 2906 -255
rect 2940 -289 2973 -255
rect 2873 -336 2973 -289
rect 3031 -255 3131 -239
rect 3031 -289 3064 -255
rect 3098 -289 3131 -255
rect 3031 -336 3131 -289
rect -3131 -583 -3031 -536
rect -3131 -617 -3098 -583
rect -3064 -617 -3031 -583
rect -3131 -633 -3031 -617
rect -2973 -583 -2873 -536
rect -2973 -617 -2940 -583
rect -2906 -617 -2873 -583
rect -2973 -633 -2873 -617
rect -2815 -583 -2715 -536
rect -2815 -617 -2782 -583
rect -2748 -617 -2715 -583
rect -2815 -633 -2715 -617
rect -2657 -583 -2557 -536
rect -2657 -617 -2624 -583
rect -2590 -617 -2557 -583
rect -2657 -633 -2557 -617
rect -2499 -583 -2399 -536
rect -2499 -617 -2466 -583
rect -2432 -617 -2399 -583
rect -2499 -633 -2399 -617
rect -2341 -583 -2241 -536
rect -2341 -617 -2308 -583
rect -2274 -617 -2241 -583
rect -2341 -633 -2241 -617
rect -2183 -583 -2083 -536
rect -2183 -617 -2150 -583
rect -2116 -617 -2083 -583
rect -2183 -633 -2083 -617
rect -2025 -583 -1925 -536
rect -2025 -617 -1992 -583
rect -1958 -617 -1925 -583
rect -2025 -633 -1925 -617
rect -1867 -583 -1767 -536
rect -1867 -617 -1834 -583
rect -1800 -617 -1767 -583
rect -1867 -633 -1767 -617
rect -1709 -583 -1609 -536
rect -1709 -617 -1676 -583
rect -1642 -617 -1609 -583
rect -1709 -633 -1609 -617
rect -1551 -583 -1451 -536
rect -1551 -617 -1518 -583
rect -1484 -617 -1451 -583
rect -1551 -633 -1451 -617
rect -1393 -583 -1293 -536
rect -1393 -617 -1360 -583
rect -1326 -617 -1293 -583
rect -1393 -633 -1293 -617
rect -1235 -583 -1135 -536
rect -1235 -617 -1202 -583
rect -1168 -617 -1135 -583
rect -1235 -633 -1135 -617
rect -1077 -583 -977 -536
rect -1077 -617 -1044 -583
rect -1010 -617 -977 -583
rect -1077 -633 -977 -617
rect -919 -583 -819 -536
rect -919 -617 -886 -583
rect -852 -617 -819 -583
rect -919 -633 -819 -617
rect -761 -583 -661 -536
rect -761 -617 -728 -583
rect -694 -617 -661 -583
rect -761 -633 -661 -617
rect -603 -583 -503 -536
rect -603 -617 -570 -583
rect -536 -617 -503 -583
rect -603 -633 -503 -617
rect -445 -583 -345 -536
rect -445 -617 -412 -583
rect -378 -617 -345 -583
rect -445 -633 -345 -617
rect -287 -583 -187 -536
rect -287 -617 -254 -583
rect -220 -617 -187 -583
rect -287 -633 -187 -617
rect -129 -583 -29 -536
rect -129 -617 -96 -583
rect -62 -617 -29 -583
rect -129 -633 -29 -617
rect 29 -583 129 -536
rect 29 -617 62 -583
rect 96 -617 129 -583
rect 29 -633 129 -617
rect 187 -583 287 -536
rect 187 -617 220 -583
rect 254 -617 287 -583
rect 187 -633 287 -617
rect 345 -583 445 -536
rect 345 -617 378 -583
rect 412 -617 445 -583
rect 345 -633 445 -617
rect 503 -583 603 -536
rect 503 -617 536 -583
rect 570 -617 603 -583
rect 503 -633 603 -617
rect 661 -583 761 -536
rect 661 -617 694 -583
rect 728 -617 761 -583
rect 661 -633 761 -617
rect 819 -583 919 -536
rect 819 -617 852 -583
rect 886 -617 919 -583
rect 819 -633 919 -617
rect 977 -583 1077 -536
rect 977 -617 1010 -583
rect 1044 -617 1077 -583
rect 977 -633 1077 -617
rect 1135 -583 1235 -536
rect 1135 -617 1168 -583
rect 1202 -617 1235 -583
rect 1135 -633 1235 -617
rect 1293 -583 1393 -536
rect 1293 -617 1326 -583
rect 1360 -617 1393 -583
rect 1293 -633 1393 -617
rect 1451 -583 1551 -536
rect 1451 -617 1484 -583
rect 1518 -617 1551 -583
rect 1451 -633 1551 -617
rect 1609 -583 1709 -536
rect 1609 -617 1642 -583
rect 1676 -617 1709 -583
rect 1609 -633 1709 -617
rect 1767 -583 1867 -536
rect 1767 -617 1800 -583
rect 1834 -617 1867 -583
rect 1767 -633 1867 -617
rect 1925 -583 2025 -536
rect 1925 -617 1958 -583
rect 1992 -617 2025 -583
rect 1925 -633 2025 -617
rect 2083 -583 2183 -536
rect 2083 -617 2116 -583
rect 2150 -617 2183 -583
rect 2083 -633 2183 -617
rect 2241 -583 2341 -536
rect 2241 -617 2274 -583
rect 2308 -617 2341 -583
rect 2241 -633 2341 -617
rect 2399 -583 2499 -536
rect 2399 -617 2432 -583
rect 2466 -617 2499 -583
rect 2399 -633 2499 -617
rect 2557 -583 2657 -536
rect 2557 -617 2590 -583
rect 2624 -617 2657 -583
rect 2557 -633 2657 -617
rect 2715 -583 2815 -536
rect 2715 -617 2748 -583
rect 2782 -617 2815 -583
rect 2715 -633 2815 -617
rect 2873 -583 2973 -536
rect 2873 -617 2906 -583
rect 2940 -617 2973 -583
rect 2873 -633 2973 -617
rect 3031 -583 3131 -536
rect 3031 -617 3064 -583
rect 3098 -617 3131 -583
rect 3031 -633 3131 -617
rect -3131 -691 -3031 -675
rect -3131 -725 -3098 -691
rect -3064 -725 -3031 -691
rect -3131 -772 -3031 -725
rect -2973 -691 -2873 -675
rect -2973 -725 -2940 -691
rect -2906 -725 -2873 -691
rect -2973 -772 -2873 -725
rect -2815 -691 -2715 -675
rect -2815 -725 -2782 -691
rect -2748 -725 -2715 -691
rect -2815 -772 -2715 -725
rect -2657 -691 -2557 -675
rect -2657 -725 -2624 -691
rect -2590 -725 -2557 -691
rect -2657 -772 -2557 -725
rect -2499 -691 -2399 -675
rect -2499 -725 -2466 -691
rect -2432 -725 -2399 -691
rect -2499 -772 -2399 -725
rect -2341 -691 -2241 -675
rect -2341 -725 -2308 -691
rect -2274 -725 -2241 -691
rect -2341 -772 -2241 -725
rect -2183 -691 -2083 -675
rect -2183 -725 -2150 -691
rect -2116 -725 -2083 -691
rect -2183 -772 -2083 -725
rect -2025 -691 -1925 -675
rect -2025 -725 -1992 -691
rect -1958 -725 -1925 -691
rect -2025 -772 -1925 -725
rect -1867 -691 -1767 -675
rect -1867 -725 -1834 -691
rect -1800 -725 -1767 -691
rect -1867 -772 -1767 -725
rect -1709 -691 -1609 -675
rect -1709 -725 -1676 -691
rect -1642 -725 -1609 -691
rect -1709 -772 -1609 -725
rect -1551 -691 -1451 -675
rect -1551 -725 -1518 -691
rect -1484 -725 -1451 -691
rect -1551 -772 -1451 -725
rect -1393 -691 -1293 -675
rect -1393 -725 -1360 -691
rect -1326 -725 -1293 -691
rect -1393 -772 -1293 -725
rect -1235 -691 -1135 -675
rect -1235 -725 -1202 -691
rect -1168 -725 -1135 -691
rect -1235 -772 -1135 -725
rect -1077 -691 -977 -675
rect -1077 -725 -1044 -691
rect -1010 -725 -977 -691
rect -1077 -772 -977 -725
rect -919 -691 -819 -675
rect -919 -725 -886 -691
rect -852 -725 -819 -691
rect -919 -772 -819 -725
rect -761 -691 -661 -675
rect -761 -725 -728 -691
rect -694 -725 -661 -691
rect -761 -772 -661 -725
rect -603 -691 -503 -675
rect -603 -725 -570 -691
rect -536 -725 -503 -691
rect -603 -772 -503 -725
rect -445 -691 -345 -675
rect -445 -725 -412 -691
rect -378 -725 -345 -691
rect -445 -772 -345 -725
rect -287 -691 -187 -675
rect -287 -725 -254 -691
rect -220 -725 -187 -691
rect -287 -772 -187 -725
rect -129 -691 -29 -675
rect -129 -725 -96 -691
rect -62 -725 -29 -691
rect -129 -772 -29 -725
rect 29 -691 129 -675
rect 29 -725 62 -691
rect 96 -725 129 -691
rect 29 -772 129 -725
rect 187 -691 287 -675
rect 187 -725 220 -691
rect 254 -725 287 -691
rect 187 -772 287 -725
rect 345 -691 445 -675
rect 345 -725 378 -691
rect 412 -725 445 -691
rect 345 -772 445 -725
rect 503 -691 603 -675
rect 503 -725 536 -691
rect 570 -725 603 -691
rect 503 -772 603 -725
rect 661 -691 761 -675
rect 661 -725 694 -691
rect 728 -725 761 -691
rect 661 -772 761 -725
rect 819 -691 919 -675
rect 819 -725 852 -691
rect 886 -725 919 -691
rect 819 -772 919 -725
rect 977 -691 1077 -675
rect 977 -725 1010 -691
rect 1044 -725 1077 -691
rect 977 -772 1077 -725
rect 1135 -691 1235 -675
rect 1135 -725 1168 -691
rect 1202 -725 1235 -691
rect 1135 -772 1235 -725
rect 1293 -691 1393 -675
rect 1293 -725 1326 -691
rect 1360 -725 1393 -691
rect 1293 -772 1393 -725
rect 1451 -691 1551 -675
rect 1451 -725 1484 -691
rect 1518 -725 1551 -691
rect 1451 -772 1551 -725
rect 1609 -691 1709 -675
rect 1609 -725 1642 -691
rect 1676 -725 1709 -691
rect 1609 -772 1709 -725
rect 1767 -691 1867 -675
rect 1767 -725 1800 -691
rect 1834 -725 1867 -691
rect 1767 -772 1867 -725
rect 1925 -691 2025 -675
rect 1925 -725 1958 -691
rect 1992 -725 2025 -691
rect 1925 -772 2025 -725
rect 2083 -691 2183 -675
rect 2083 -725 2116 -691
rect 2150 -725 2183 -691
rect 2083 -772 2183 -725
rect 2241 -691 2341 -675
rect 2241 -725 2274 -691
rect 2308 -725 2341 -691
rect 2241 -772 2341 -725
rect 2399 -691 2499 -675
rect 2399 -725 2432 -691
rect 2466 -725 2499 -691
rect 2399 -772 2499 -725
rect 2557 -691 2657 -675
rect 2557 -725 2590 -691
rect 2624 -725 2657 -691
rect 2557 -772 2657 -725
rect 2715 -691 2815 -675
rect 2715 -725 2748 -691
rect 2782 -725 2815 -691
rect 2715 -772 2815 -725
rect 2873 -691 2973 -675
rect 2873 -725 2906 -691
rect 2940 -725 2973 -691
rect 2873 -772 2973 -725
rect 3031 -691 3131 -675
rect 3031 -725 3064 -691
rect 3098 -725 3131 -691
rect 3031 -772 3131 -725
rect -3131 -1019 -3031 -972
rect -3131 -1053 -3098 -1019
rect -3064 -1053 -3031 -1019
rect -3131 -1069 -3031 -1053
rect -2973 -1019 -2873 -972
rect -2973 -1053 -2940 -1019
rect -2906 -1053 -2873 -1019
rect -2973 -1069 -2873 -1053
rect -2815 -1019 -2715 -972
rect -2815 -1053 -2782 -1019
rect -2748 -1053 -2715 -1019
rect -2815 -1069 -2715 -1053
rect -2657 -1019 -2557 -972
rect -2657 -1053 -2624 -1019
rect -2590 -1053 -2557 -1019
rect -2657 -1069 -2557 -1053
rect -2499 -1019 -2399 -972
rect -2499 -1053 -2466 -1019
rect -2432 -1053 -2399 -1019
rect -2499 -1069 -2399 -1053
rect -2341 -1019 -2241 -972
rect -2341 -1053 -2308 -1019
rect -2274 -1053 -2241 -1019
rect -2341 -1069 -2241 -1053
rect -2183 -1019 -2083 -972
rect -2183 -1053 -2150 -1019
rect -2116 -1053 -2083 -1019
rect -2183 -1069 -2083 -1053
rect -2025 -1019 -1925 -972
rect -2025 -1053 -1992 -1019
rect -1958 -1053 -1925 -1019
rect -2025 -1069 -1925 -1053
rect -1867 -1019 -1767 -972
rect -1867 -1053 -1834 -1019
rect -1800 -1053 -1767 -1019
rect -1867 -1069 -1767 -1053
rect -1709 -1019 -1609 -972
rect -1709 -1053 -1676 -1019
rect -1642 -1053 -1609 -1019
rect -1709 -1069 -1609 -1053
rect -1551 -1019 -1451 -972
rect -1551 -1053 -1518 -1019
rect -1484 -1053 -1451 -1019
rect -1551 -1069 -1451 -1053
rect -1393 -1019 -1293 -972
rect -1393 -1053 -1360 -1019
rect -1326 -1053 -1293 -1019
rect -1393 -1069 -1293 -1053
rect -1235 -1019 -1135 -972
rect -1235 -1053 -1202 -1019
rect -1168 -1053 -1135 -1019
rect -1235 -1069 -1135 -1053
rect -1077 -1019 -977 -972
rect -1077 -1053 -1044 -1019
rect -1010 -1053 -977 -1019
rect -1077 -1069 -977 -1053
rect -919 -1019 -819 -972
rect -919 -1053 -886 -1019
rect -852 -1053 -819 -1019
rect -919 -1069 -819 -1053
rect -761 -1019 -661 -972
rect -761 -1053 -728 -1019
rect -694 -1053 -661 -1019
rect -761 -1069 -661 -1053
rect -603 -1019 -503 -972
rect -603 -1053 -570 -1019
rect -536 -1053 -503 -1019
rect -603 -1069 -503 -1053
rect -445 -1019 -345 -972
rect -445 -1053 -412 -1019
rect -378 -1053 -345 -1019
rect -445 -1069 -345 -1053
rect -287 -1019 -187 -972
rect -287 -1053 -254 -1019
rect -220 -1053 -187 -1019
rect -287 -1069 -187 -1053
rect -129 -1019 -29 -972
rect -129 -1053 -96 -1019
rect -62 -1053 -29 -1019
rect -129 -1069 -29 -1053
rect 29 -1019 129 -972
rect 29 -1053 62 -1019
rect 96 -1053 129 -1019
rect 29 -1069 129 -1053
rect 187 -1019 287 -972
rect 187 -1053 220 -1019
rect 254 -1053 287 -1019
rect 187 -1069 287 -1053
rect 345 -1019 445 -972
rect 345 -1053 378 -1019
rect 412 -1053 445 -1019
rect 345 -1069 445 -1053
rect 503 -1019 603 -972
rect 503 -1053 536 -1019
rect 570 -1053 603 -1019
rect 503 -1069 603 -1053
rect 661 -1019 761 -972
rect 661 -1053 694 -1019
rect 728 -1053 761 -1019
rect 661 -1069 761 -1053
rect 819 -1019 919 -972
rect 819 -1053 852 -1019
rect 886 -1053 919 -1019
rect 819 -1069 919 -1053
rect 977 -1019 1077 -972
rect 977 -1053 1010 -1019
rect 1044 -1053 1077 -1019
rect 977 -1069 1077 -1053
rect 1135 -1019 1235 -972
rect 1135 -1053 1168 -1019
rect 1202 -1053 1235 -1019
rect 1135 -1069 1235 -1053
rect 1293 -1019 1393 -972
rect 1293 -1053 1326 -1019
rect 1360 -1053 1393 -1019
rect 1293 -1069 1393 -1053
rect 1451 -1019 1551 -972
rect 1451 -1053 1484 -1019
rect 1518 -1053 1551 -1019
rect 1451 -1069 1551 -1053
rect 1609 -1019 1709 -972
rect 1609 -1053 1642 -1019
rect 1676 -1053 1709 -1019
rect 1609 -1069 1709 -1053
rect 1767 -1019 1867 -972
rect 1767 -1053 1800 -1019
rect 1834 -1053 1867 -1019
rect 1767 -1069 1867 -1053
rect 1925 -1019 2025 -972
rect 1925 -1053 1958 -1019
rect 1992 -1053 2025 -1019
rect 1925 -1069 2025 -1053
rect 2083 -1019 2183 -972
rect 2083 -1053 2116 -1019
rect 2150 -1053 2183 -1019
rect 2083 -1069 2183 -1053
rect 2241 -1019 2341 -972
rect 2241 -1053 2274 -1019
rect 2308 -1053 2341 -1019
rect 2241 -1069 2341 -1053
rect 2399 -1019 2499 -972
rect 2399 -1053 2432 -1019
rect 2466 -1053 2499 -1019
rect 2399 -1069 2499 -1053
rect 2557 -1019 2657 -972
rect 2557 -1053 2590 -1019
rect 2624 -1053 2657 -1019
rect 2557 -1069 2657 -1053
rect 2715 -1019 2815 -972
rect 2715 -1053 2748 -1019
rect 2782 -1053 2815 -1019
rect 2715 -1069 2815 -1053
rect 2873 -1019 2973 -972
rect 2873 -1053 2906 -1019
rect 2940 -1053 2973 -1019
rect 2873 -1069 2973 -1053
rect 3031 -1019 3131 -972
rect 3031 -1053 3064 -1019
rect 3098 -1053 3131 -1019
rect 3031 -1069 3131 -1053
<< polycont >>
rect -3098 1019 -3064 1053
rect -2940 1019 -2906 1053
rect -2782 1019 -2748 1053
rect -2624 1019 -2590 1053
rect -2466 1019 -2432 1053
rect -2308 1019 -2274 1053
rect -2150 1019 -2116 1053
rect -1992 1019 -1958 1053
rect -1834 1019 -1800 1053
rect -1676 1019 -1642 1053
rect -1518 1019 -1484 1053
rect -1360 1019 -1326 1053
rect -1202 1019 -1168 1053
rect -1044 1019 -1010 1053
rect -886 1019 -852 1053
rect -728 1019 -694 1053
rect -570 1019 -536 1053
rect -412 1019 -378 1053
rect -254 1019 -220 1053
rect -96 1019 -62 1053
rect 62 1019 96 1053
rect 220 1019 254 1053
rect 378 1019 412 1053
rect 536 1019 570 1053
rect 694 1019 728 1053
rect 852 1019 886 1053
rect 1010 1019 1044 1053
rect 1168 1019 1202 1053
rect 1326 1019 1360 1053
rect 1484 1019 1518 1053
rect 1642 1019 1676 1053
rect 1800 1019 1834 1053
rect 1958 1019 1992 1053
rect 2116 1019 2150 1053
rect 2274 1019 2308 1053
rect 2432 1019 2466 1053
rect 2590 1019 2624 1053
rect 2748 1019 2782 1053
rect 2906 1019 2940 1053
rect 3064 1019 3098 1053
rect -3098 691 -3064 725
rect -2940 691 -2906 725
rect -2782 691 -2748 725
rect -2624 691 -2590 725
rect -2466 691 -2432 725
rect -2308 691 -2274 725
rect -2150 691 -2116 725
rect -1992 691 -1958 725
rect -1834 691 -1800 725
rect -1676 691 -1642 725
rect -1518 691 -1484 725
rect -1360 691 -1326 725
rect -1202 691 -1168 725
rect -1044 691 -1010 725
rect -886 691 -852 725
rect -728 691 -694 725
rect -570 691 -536 725
rect -412 691 -378 725
rect -254 691 -220 725
rect -96 691 -62 725
rect 62 691 96 725
rect 220 691 254 725
rect 378 691 412 725
rect 536 691 570 725
rect 694 691 728 725
rect 852 691 886 725
rect 1010 691 1044 725
rect 1168 691 1202 725
rect 1326 691 1360 725
rect 1484 691 1518 725
rect 1642 691 1676 725
rect 1800 691 1834 725
rect 1958 691 1992 725
rect 2116 691 2150 725
rect 2274 691 2308 725
rect 2432 691 2466 725
rect 2590 691 2624 725
rect 2748 691 2782 725
rect 2906 691 2940 725
rect 3064 691 3098 725
rect -3098 583 -3064 617
rect -2940 583 -2906 617
rect -2782 583 -2748 617
rect -2624 583 -2590 617
rect -2466 583 -2432 617
rect -2308 583 -2274 617
rect -2150 583 -2116 617
rect -1992 583 -1958 617
rect -1834 583 -1800 617
rect -1676 583 -1642 617
rect -1518 583 -1484 617
rect -1360 583 -1326 617
rect -1202 583 -1168 617
rect -1044 583 -1010 617
rect -886 583 -852 617
rect -728 583 -694 617
rect -570 583 -536 617
rect -412 583 -378 617
rect -254 583 -220 617
rect -96 583 -62 617
rect 62 583 96 617
rect 220 583 254 617
rect 378 583 412 617
rect 536 583 570 617
rect 694 583 728 617
rect 852 583 886 617
rect 1010 583 1044 617
rect 1168 583 1202 617
rect 1326 583 1360 617
rect 1484 583 1518 617
rect 1642 583 1676 617
rect 1800 583 1834 617
rect 1958 583 1992 617
rect 2116 583 2150 617
rect 2274 583 2308 617
rect 2432 583 2466 617
rect 2590 583 2624 617
rect 2748 583 2782 617
rect 2906 583 2940 617
rect 3064 583 3098 617
rect -3098 255 -3064 289
rect -2940 255 -2906 289
rect -2782 255 -2748 289
rect -2624 255 -2590 289
rect -2466 255 -2432 289
rect -2308 255 -2274 289
rect -2150 255 -2116 289
rect -1992 255 -1958 289
rect -1834 255 -1800 289
rect -1676 255 -1642 289
rect -1518 255 -1484 289
rect -1360 255 -1326 289
rect -1202 255 -1168 289
rect -1044 255 -1010 289
rect -886 255 -852 289
rect -728 255 -694 289
rect -570 255 -536 289
rect -412 255 -378 289
rect -254 255 -220 289
rect -96 255 -62 289
rect 62 255 96 289
rect 220 255 254 289
rect 378 255 412 289
rect 536 255 570 289
rect 694 255 728 289
rect 852 255 886 289
rect 1010 255 1044 289
rect 1168 255 1202 289
rect 1326 255 1360 289
rect 1484 255 1518 289
rect 1642 255 1676 289
rect 1800 255 1834 289
rect 1958 255 1992 289
rect 2116 255 2150 289
rect 2274 255 2308 289
rect 2432 255 2466 289
rect 2590 255 2624 289
rect 2748 255 2782 289
rect 2906 255 2940 289
rect 3064 255 3098 289
rect -3098 147 -3064 181
rect -2940 147 -2906 181
rect -2782 147 -2748 181
rect -2624 147 -2590 181
rect -2466 147 -2432 181
rect -2308 147 -2274 181
rect -2150 147 -2116 181
rect -1992 147 -1958 181
rect -1834 147 -1800 181
rect -1676 147 -1642 181
rect -1518 147 -1484 181
rect -1360 147 -1326 181
rect -1202 147 -1168 181
rect -1044 147 -1010 181
rect -886 147 -852 181
rect -728 147 -694 181
rect -570 147 -536 181
rect -412 147 -378 181
rect -254 147 -220 181
rect -96 147 -62 181
rect 62 147 96 181
rect 220 147 254 181
rect 378 147 412 181
rect 536 147 570 181
rect 694 147 728 181
rect 852 147 886 181
rect 1010 147 1044 181
rect 1168 147 1202 181
rect 1326 147 1360 181
rect 1484 147 1518 181
rect 1642 147 1676 181
rect 1800 147 1834 181
rect 1958 147 1992 181
rect 2116 147 2150 181
rect 2274 147 2308 181
rect 2432 147 2466 181
rect 2590 147 2624 181
rect 2748 147 2782 181
rect 2906 147 2940 181
rect 3064 147 3098 181
rect -3098 -181 -3064 -147
rect -2940 -181 -2906 -147
rect -2782 -181 -2748 -147
rect -2624 -181 -2590 -147
rect -2466 -181 -2432 -147
rect -2308 -181 -2274 -147
rect -2150 -181 -2116 -147
rect -1992 -181 -1958 -147
rect -1834 -181 -1800 -147
rect -1676 -181 -1642 -147
rect -1518 -181 -1484 -147
rect -1360 -181 -1326 -147
rect -1202 -181 -1168 -147
rect -1044 -181 -1010 -147
rect -886 -181 -852 -147
rect -728 -181 -694 -147
rect -570 -181 -536 -147
rect -412 -181 -378 -147
rect -254 -181 -220 -147
rect -96 -181 -62 -147
rect 62 -181 96 -147
rect 220 -181 254 -147
rect 378 -181 412 -147
rect 536 -181 570 -147
rect 694 -181 728 -147
rect 852 -181 886 -147
rect 1010 -181 1044 -147
rect 1168 -181 1202 -147
rect 1326 -181 1360 -147
rect 1484 -181 1518 -147
rect 1642 -181 1676 -147
rect 1800 -181 1834 -147
rect 1958 -181 1992 -147
rect 2116 -181 2150 -147
rect 2274 -181 2308 -147
rect 2432 -181 2466 -147
rect 2590 -181 2624 -147
rect 2748 -181 2782 -147
rect 2906 -181 2940 -147
rect 3064 -181 3098 -147
rect -3098 -289 -3064 -255
rect -2940 -289 -2906 -255
rect -2782 -289 -2748 -255
rect -2624 -289 -2590 -255
rect -2466 -289 -2432 -255
rect -2308 -289 -2274 -255
rect -2150 -289 -2116 -255
rect -1992 -289 -1958 -255
rect -1834 -289 -1800 -255
rect -1676 -289 -1642 -255
rect -1518 -289 -1484 -255
rect -1360 -289 -1326 -255
rect -1202 -289 -1168 -255
rect -1044 -289 -1010 -255
rect -886 -289 -852 -255
rect -728 -289 -694 -255
rect -570 -289 -536 -255
rect -412 -289 -378 -255
rect -254 -289 -220 -255
rect -96 -289 -62 -255
rect 62 -289 96 -255
rect 220 -289 254 -255
rect 378 -289 412 -255
rect 536 -289 570 -255
rect 694 -289 728 -255
rect 852 -289 886 -255
rect 1010 -289 1044 -255
rect 1168 -289 1202 -255
rect 1326 -289 1360 -255
rect 1484 -289 1518 -255
rect 1642 -289 1676 -255
rect 1800 -289 1834 -255
rect 1958 -289 1992 -255
rect 2116 -289 2150 -255
rect 2274 -289 2308 -255
rect 2432 -289 2466 -255
rect 2590 -289 2624 -255
rect 2748 -289 2782 -255
rect 2906 -289 2940 -255
rect 3064 -289 3098 -255
rect -3098 -617 -3064 -583
rect -2940 -617 -2906 -583
rect -2782 -617 -2748 -583
rect -2624 -617 -2590 -583
rect -2466 -617 -2432 -583
rect -2308 -617 -2274 -583
rect -2150 -617 -2116 -583
rect -1992 -617 -1958 -583
rect -1834 -617 -1800 -583
rect -1676 -617 -1642 -583
rect -1518 -617 -1484 -583
rect -1360 -617 -1326 -583
rect -1202 -617 -1168 -583
rect -1044 -617 -1010 -583
rect -886 -617 -852 -583
rect -728 -617 -694 -583
rect -570 -617 -536 -583
rect -412 -617 -378 -583
rect -254 -617 -220 -583
rect -96 -617 -62 -583
rect 62 -617 96 -583
rect 220 -617 254 -583
rect 378 -617 412 -583
rect 536 -617 570 -583
rect 694 -617 728 -583
rect 852 -617 886 -583
rect 1010 -617 1044 -583
rect 1168 -617 1202 -583
rect 1326 -617 1360 -583
rect 1484 -617 1518 -583
rect 1642 -617 1676 -583
rect 1800 -617 1834 -583
rect 1958 -617 1992 -583
rect 2116 -617 2150 -583
rect 2274 -617 2308 -583
rect 2432 -617 2466 -583
rect 2590 -617 2624 -583
rect 2748 -617 2782 -583
rect 2906 -617 2940 -583
rect 3064 -617 3098 -583
rect -3098 -725 -3064 -691
rect -2940 -725 -2906 -691
rect -2782 -725 -2748 -691
rect -2624 -725 -2590 -691
rect -2466 -725 -2432 -691
rect -2308 -725 -2274 -691
rect -2150 -725 -2116 -691
rect -1992 -725 -1958 -691
rect -1834 -725 -1800 -691
rect -1676 -725 -1642 -691
rect -1518 -725 -1484 -691
rect -1360 -725 -1326 -691
rect -1202 -725 -1168 -691
rect -1044 -725 -1010 -691
rect -886 -725 -852 -691
rect -728 -725 -694 -691
rect -570 -725 -536 -691
rect -412 -725 -378 -691
rect -254 -725 -220 -691
rect -96 -725 -62 -691
rect 62 -725 96 -691
rect 220 -725 254 -691
rect 378 -725 412 -691
rect 536 -725 570 -691
rect 694 -725 728 -691
rect 852 -725 886 -691
rect 1010 -725 1044 -691
rect 1168 -725 1202 -691
rect 1326 -725 1360 -691
rect 1484 -725 1518 -691
rect 1642 -725 1676 -691
rect 1800 -725 1834 -691
rect 1958 -725 1992 -691
rect 2116 -725 2150 -691
rect 2274 -725 2308 -691
rect 2432 -725 2466 -691
rect 2590 -725 2624 -691
rect 2748 -725 2782 -691
rect 2906 -725 2940 -691
rect 3064 -725 3098 -691
rect -3098 -1053 -3064 -1019
rect -2940 -1053 -2906 -1019
rect -2782 -1053 -2748 -1019
rect -2624 -1053 -2590 -1019
rect -2466 -1053 -2432 -1019
rect -2308 -1053 -2274 -1019
rect -2150 -1053 -2116 -1019
rect -1992 -1053 -1958 -1019
rect -1834 -1053 -1800 -1019
rect -1676 -1053 -1642 -1019
rect -1518 -1053 -1484 -1019
rect -1360 -1053 -1326 -1019
rect -1202 -1053 -1168 -1019
rect -1044 -1053 -1010 -1019
rect -886 -1053 -852 -1019
rect -728 -1053 -694 -1019
rect -570 -1053 -536 -1019
rect -412 -1053 -378 -1019
rect -254 -1053 -220 -1019
rect -96 -1053 -62 -1019
rect 62 -1053 96 -1019
rect 220 -1053 254 -1019
rect 378 -1053 412 -1019
rect 536 -1053 570 -1019
rect 694 -1053 728 -1019
rect 852 -1053 886 -1019
rect 1010 -1053 1044 -1019
rect 1168 -1053 1202 -1019
rect 1326 -1053 1360 -1019
rect 1484 -1053 1518 -1019
rect 1642 -1053 1676 -1019
rect 1800 -1053 1834 -1019
rect 1958 -1053 1992 -1019
rect 2116 -1053 2150 -1019
rect 2274 -1053 2308 -1019
rect 2432 -1053 2466 -1019
rect 2590 -1053 2624 -1019
rect 2748 -1053 2782 -1019
rect 2906 -1053 2940 -1019
rect 3064 -1053 3098 -1019
<< locali >>
rect -3311 1157 -3213 1191
rect -3179 1157 -3145 1191
rect -3111 1157 -3077 1191
rect -3043 1157 -3009 1191
rect -2975 1157 -2941 1191
rect -2907 1157 -2873 1191
rect -2839 1157 -2805 1191
rect -2771 1157 -2737 1191
rect -2703 1157 -2669 1191
rect -2635 1157 -2601 1191
rect -2567 1157 -2533 1191
rect -2499 1157 -2465 1191
rect -2431 1157 -2397 1191
rect -2363 1157 -2329 1191
rect -2295 1157 -2261 1191
rect -2227 1157 -2193 1191
rect -2159 1157 -2125 1191
rect -2091 1157 -2057 1191
rect -2023 1157 -1989 1191
rect -1955 1157 -1921 1191
rect -1887 1157 -1853 1191
rect -1819 1157 -1785 1191
rect -1751 1157 -1717 1191
rect -1683 1157 -1649 1191
rect -1615 1157 -1581 1191
rect -1547 1157 -1513 1191
rect -1479 1157 -1445 1191
rect -1411 1157 -1377 1191
rect -1343 1157 -1309 1191
rect -1275 1157 -1241 1191
rect -1207 1157 -1173 1191
rect -1139 1157 -1105 1191
rect -1071 1157 -1037 1191
rect -1003 1157 -969 1191
rect -935 1157 -901 1191
rect -867 1157 -833 1191
rect -799 1157 -765 1191
rect -731 1157 -697 1191
rect -663 1157 -629 1191
rect -595 1157 -561 1191
rect -527 1157 -493 1191
rect -459 1157 -425 1191
rect -391 1157 -357 1191
rect -323 1157 -289 1191
rect -255 1157 -221 1191
rect -187 1157 -153 1191
rect -119 1157 -85 1191
rect -51 1157 -17 1191
rect 17 1157 51 1191
rect 85 1157 119 1191
rect 153 1157 187 1191
rect 221 1157 255 1191
rect 289 1157 323 1191
rect 357 1157 391 1191
rect 425 1157 459 1191
rect 493 1157 527 1191
rect 561 1157 595 1191
rect 629 1157 663 1191
rect 697 1157 731 1191
rect 765 1157 799 1191
rect 833 1157 867 1191
rect 901 1157 935 1191
rect 969 1157 1003 1191
rect 1037 1157 1071 1191
rect 1105 1157 1139 1191
rect 1173 1157 1207 1191
rect 1241 1157 1275 1191
rect 1309 1157 1343 1191
rect 1377 1157 1411 1191
rect 1445 1157 1479 1191
rect 1513 1157 1547 1191
rect 1581 1157 1615 1191
rect 1649 1157 1683 1191
rect 1717 1157 1751 1191
rect 1785 1157 1819 1191
rect 1853 1157 1887 1191
rect 1921 1157 1955 1191
rect 1989 1157 2023 1191
rect 2057 1157 2091 1191
rect 2125 1157 2159 1191
rect 2193 1157 2227 1191
rect 2261 1157 2295 1191
rect 2329 1157 2363 1191
rect 2397 1157 2431 1191
rect 2465 1157 2499 1191
rect 2533 1157 2567 1191
rect 2601 1157 2635 1191
rect 2669 1157 2703 1191
rect 2737 1157 2771 1191
rect 2805 1157 2839 1191
rect 2873 1157 2907 1191
rect 2941 1157 2975 1191
rect 3009 1157 3043 1191
rect 3077 1157 3111 1191
rect 3145 1157 3179 1191
rect 3213 1157 3311 1191
rect -3311 1071 -3277 1157
rect 3277 1071 3311 1157
rect -3311 1003 -3277 1037
rect -3131 1019 -3098 1053
rect -3064 1019 -3031 1053
rect -2973 1019 -2940 1053
rect -2906 1019 -2873 1053
rect -2815 1019 -2782 1053
rect -2748 1019 -2715 1053
rect -2657 1019 -2624 1053
rect -2590 1019 -2557 1053
rect -2499 1019 -2466 1053
rect -2432 1019 -2399 1053
rect -2341 1019 -2308 1053
rect -2274 1019 -2241 1053
rect -2183 1019 -2150 1053
rect -2116 1019 -2083 1053
rect -2025 1019 -1992 1053
rect -1958 1019 -1925 1053
rect -1867 1019 -1834 1053
rect -1800 1019 -1767 1053
rect -1709 1019 -1676 1053
rect -1642 1019 -1609 1053
rect -1551 1019 -1518 1053
rect -1484 1019 -1451 1053
rect -1393 1019 -1360 1053
rect -1326 1019 -1293 1053
rect -1235 1019 -1202 1053
rect -1168 1019 -1135 1053
rect -1077 1019 -1044 1053
rect -1010 1019 -977 1053
rect -919 1019 -886 1053
rect -852 1019 -819 1053
rect -761 1019 -728 1053
rect -694 1019 -661 1053
rect -603 1019 -570 1053
rect -536 1019 -503 1053
rect -445 1019 -412 1053
rect -378 1019 -345 1053
rect -287 1019 -254 1053
rect -220 1019 -187 1053
rect -129 1019 -96 1053
rect -62 1019 -29 1053
rect 29 1019 62 1053
rect 96 1019 129 1053
rect 187 1019 220 1053
rect 254 1019 287 1053
rect 345 1019 378 1053
rect 412 1019 445 1053
rect 503 1019 536 1053
rect 570 1019 603 1053
rect 661 1019 694 1053
rect 728 1019 761 1053
rect 819 1019 852 1053
rect 886 1019 919 1053
rect 977 1019 1010 1053
rect 1044 1019 1077 1053
rect 1135 1019 1168 1053
rect 1202 1019 1235 1053
rect 1293 1019 1326 1053
rect 1360 1019 1393 1053
rect 1451 1019 1484 1053
rect 1518 1019 1551 1053
rect 1609 1019 1642 1053
rect 1676 1019 1709 1053
rect 1767 1019 1800 1053
rect 1834 1019 1867 1053
rect 1925 1019 1958 1053
rect 1992 1019 2025 1053
rect 2083 1019 2116 1053
rect 2150 1019 2183 1053
rect 2241 1019 2274 1053
rect 2308 1019 2341 1053
rect 2399 1019 2432 1053
rect 2466 1019 2499 1053
rect 2557 1019 2590 1053
rect 2624 1019 2657 1053
rect 2715 1019 2748 1053
rect 2782 1019 2815 1053
rect 2873 1019 2906 1053
rect 2940 1019 2973 1053
rect 3031 1019 3064 1053
rect 3098 1019 3131 1053
rect 3277 1003 3311 1037
rect -3311 935 -3277 969
rect -3311 867 -3277 901
rect -3311 799 -3277 833
rect -3177 957 -3143 976
rect -3177 889 -3143 891
rect -3177 853 -3143 855
rect -3177 768 -3143 787
rect -3019 957 -2985 976
rect -3019 889 -2985 891
rect -3019 853 -2985 855
rect -3019 768 -2985 787
rect -2861 957 -2827 976
rect -2861 889 -2827 891
rect -2861 853 -2827 855
rect -2861 768 -2827 787
rect -2703 957 -2669 976
rect -2703 889 -2669 891
rect -2703 853 -2669 855
rect -2703 768 -2669 787
rect -2545 957 -2511 976
rect -2545 889 -2511 891
rect -2545 853 -2511 855
rect -2545 768 -2511 787
rect -2387 957 -2353 976
rect -2387 889 -2353 891
rect -2387 853 -2353 855
rect -2387 768 -2353 787
rect -2229 957 -2195 976
rect -2229 889 -2195 891
rect -2229 853 -2195 855
rect -2229 768 -2195 787
rect -2071 957 -2037 976
rect -2071 889 -2037 891
rect -2071 853 -2037 855
rect -2071 768 -2037 787
rect -1913 957 -1879 976
rect -1913 889 -1879 891
rect -1913 853 -1879 855
rect -1913 768 -1879 787
rect -1755 957 -1721 976
rect -1755 889 -1721 891
rect -1755 853 -1721 855
rect -1755 768 -1721 787
rect -1597 957 -1563 976
rect -1597 889 -1563 891
rect -1597 853 -1563 855
rect -1597 768 -1563 787
rect -1439 957 -1405 976
rect -1439 889 -1405 891
rect -1439 853 -1405 855
rect -1439 768 -1405 787
rect -1281 957 -1247 976
rect -1281 889 -1247 891
rect -1281 853 -1247 855
rect -1281 768 -1247 787
rect -1123 957 -1089 976
rect -1123 889 -1089 891
rect -1123 853 -1089 855
rect -1123 768 -1089 787
rect -965 957 -931 976
rect -965 889 -931 891
rect -965 853 -931 855
rect -965 768 -931 787
rect -807 957 -773 976
rect -807 889 -773 891
rect -807 853 -773 855
rect -807 768 -773 787
rect -649 957 -615 976
rect -649 889 -615 891
rect -649 853 -615 855
rect -649 768 -615 787
rect -491 957 -457 976
rect -491 889 -457 891
rect -491 853 -457 855
rect -491 768 -457 787
rect -333 957 -299 976
rect -333 889 -299 891
rect -333 853 -299 855
rect -333 768 -299 787
rect -175 957 -141 976
rect -175 889 -141 891
rect -175 853 -141 855
rect -175 768 -141 787
rect -17 957 17 976
rect -17 889 17 891
rect -17 853 17 855
rect -17 768 17 787
rect 141 957 175 976
rect 141 889 175 891
rect 141 853 175 855
rect 141 768 175 787
rect 299 957 333 976
rect 299 889 333 891
rect 299 853 333 855
rect 299 768 333 787
rect 457 957 491 976
rect 457 889 491 891
rect 457 853 491 855
rect 457 768 491 787
rect 615 957 649 976
rect 615 889 649 891
rect 615 853 649 855
rect 615 768 649 787
rect 773 957 807 976
rect 773 889 807 891
rect 773 853 807 855
rect 773 768 807 787
rect 931 957 965 976
rect 931 889 965 891
rect 931 853 965 855
rect 931 768 965 787
rect 1089 957 1123 976
rect 1089 889 1123 891
rect 1089 853 1123 855
rect 1089 768 1123 787
rect 1247 957 1281 976
rect 1247 889 1281 891
rect 1247 853 1281 855
rect 1247 768 1281 787
rect 1405 957 1439 976
rect 1405 889 1439 891
rect 1405 853 1439 855
rect 1405 768 1439 787
rect 1563 957 1597 976
rect 1563 889 1597 891
rect 1563 853 1597 855
rect 1563 768 1597 787
rect 1721 957 1755 976
rect 1721 889 1755 891
rect 1721 853 1755 855
rect 1721 768 1755 787
rect 1879 957 1913 976
rect 1879 889 1913 891
rect 1879 853 1913 855
rect 1879 768 1913 787
rect 2037 957 2071 976
rect 2037 889 2071 891
rect 2037 853 2071 855
rect 2037 768 2071 787
rect 2195 957 2229 976
rect 2195 889 2229 891
rect 2195 853 2229 855
rect 2195 768 2229 787
rect 2353 957 2387 976
rect 2353 889 2387 891
rect 2353 853 2387 855
rect 2353 768 2387 787
rect 2511 957 2545 976
rect 2511 889 2545 891
rect 2511 853 2545 855
rect 2511 768 2545 787
rect 2669 957 2703 976
rect 2669 889 2703 891
rect 2669 853 2703 855
rect 2669 768 2703 787
rect 2827 957 2861 976
rect 2827 889 2861 891
rect 2827 853 2861 855
rect 2827 768 2861 787
rect 2985 957 3019 976
rect 2985 889 3019 891
rect 2985 853 3019 855
rect 2985 768 3019 787
rect 3143 957 3177 976
rect 3143 889 3177 891
rect 3143 853 3177 855
rect 3143 768 3177 787
rect 3277 935 3311 969
rect 3277 867 3311 901
rect 3277 799 3311 833
rect -3311 731 -3277 765
rect 3277 731 3311 765
rect -3311 663 -3277 697
rect -3131 691 -3098 725
rect -3064 691 -3031 725
rect -2973 691 -2940 725
rect -2906 691 -2873 725
rect -2815 691 -2782 725
rect -2748 691 -2715 725
rect -2657 691 -2624 725
rect -2590 691 -2557 725
rect -2499 691 -2466 725
rect -2432 691 -2399 725
rect -2341 691 -2308 725
rect -2274 691 -2241 725
rect -2183 691 -2150 725
rect -2116 691 -2083 725
rect -2025 691 -1992 725
rect -1958 691 -1925 725
rect -1867 691 -1834 725
rect -1800 691 -1767 725
rect -1709 691 -1676 725
rect -1642 691 -1609 725
rect -1551 691 -1518 725
rect -1484 691 -1451 725
rect -1393 691 -1360 725
rect -1326 691 -1293 725
rect -1235 691 -1202 725
rect -1168 691 -1135 725
rect -1077 691 -1044 725
rect -1010 691 -977 725
rect -919 691 -886 725
rect -852 691 -819 725
rect -761 691 -728 725
rect -694 691 -661 725
rect -603 691 -570 725
rect -536 691 -503 725
rect -445 691 -412 725
rect -378 691 -345 725
rect -287 691 -254 725
rect -220 691 -187 725
rect -129 691 -96 725
rect -62 691 -29 725
rect 29 691 62 725
rect 96 691 129 725
rect 187 691 220 725
rect 254 691 287 725
rect 345 691 378 725
rect 412 691 445 725
rect 503 691 536 725
rect 570 691 603 725
rect 661 691 694 725
rect 728 691 761 725
rect 819 691 852 725
rect 886 691 919 725
rect 977 691 1010 725
rect 1044 691 1077 725
rect 1135 691 1168 725
rect 1202 691 1235 725
rect 1293 691 1326 725
rect 1360 691 1393 725
rect 1451 691 1484 725
rect 1518 691 1551 725
rect 1609 691 1642 725
rect 1676 691 1709 725
rect 1767 691 1800 725
rect 1834 691 1867 725
rect 1925 691 1958 725
rect 1992 691 2025 725
rect 2083 691 2116 725
rect 2150 691 2183 725
rect 2241 691 2274 725
rect 2308 691 2341 725
rect 2399 691 2432 725
rect 2466 691 2499 725
rect 2557 691 2590 725
rect 2624 691 2657 725
rect 2715 691 2748 725
rect 2782 691 2815 725
rect 2873 691 2906 725
rect 2940 691 2973 725
rect 3031 691 3064 725
rect 3098 691 3131 725
rect -3311 595 -3277 629
rect 3277 663 3311 697
rect -3131 583 -3098 617
rect -3064 583 -3031 617
rect -2973 583 -2940 617
rect -2906 583 -2873 617
rect -2815 583 -2782 617
rect -2748 583 -2715 617
rect -2657 583 -2624 617
rect -2590 583 -2557 617
rect -2499 583 -2466 617
rect -2432 583 -2399 617
rect -2341 583 -2308 617
rect -2274 583 -2241 617
rect -2183 583 -2150 617
rect -2116 583 -2083 617
rect -2025 583 -1992 617
rect -1958 583 -1925 617
rect -1867 583 -1834 617
rect -1800 583 -1767 617
rect -1709 583 -1676 617
rect -1642 583 -1609 617
rect -1551 583 -1518 617
rect -1484 583 -1451 617
rect -1393 583 -1360 617
rect -1326 583 -1293 617
rect -1235 583 -1202 617
rect -1168 583 -1135 617
rect -1077 583 -1044 617
rect -1010 583 -977 617
rect -919 583 -886 617
rect -852 583 -819 617
rect -761 583 -728 617
rect -694 583 -661 617
rect -603 583 -570 617
rect -536 583 -503 617
rect -445 583 -412 617
rect -378 583 -345 617
rect -287 583 -254 617
rect -220 583 -187 617
rect -129 583 -96 617
rect -62 583 -29 617
rect 29 583 62 617
rect 96 583 129 617
rect 187 583 220 617
rect 254 583 287 617
rect 345 583 378 617
rect 412 583 445 617
rect 503 583 536 617
rect 570 583 603 617
rect 661 583 694 617
rect 728 583 761 617
rect 819 583 852 617
rect 886 583 919 617
rect 977 583 1010 617
rect 1044 583 1077 617
rect 1135 583 1168 617
rect 1202 583 1235 617
rect 1293 583 1326 617
rect 1360 583 1393 617
rect 1451 583 1484 617
rect 1518 583 1551 617
rect 1609 583 1642 617
rect 1676 583 1709 617
rect 1767 583 1800 617
rect 1834 583 1867 617
rect 1925 583 1958 617
rect 1992 583 2025 617
rect 2083 583 2116 617
rect 2150 583 2183 617
rect 2241 583 2274 617
rect 2308 583 2341 617
rect 2399 583 2432 617
rect 2466 583 2499 617
rect 2557 583 2590 617
rect 2624 583 2657 617
rect 2715 583 2748 617
rect 2782 583 2815 617
rect 2873 583 2906 617
rect 2940 583 2973 617
rect 3031 583 3064 617
rect 3098 583 3131 617
rect 3277 595 3311 629
rect -3311 527 -3277 561
rect -3311 459 -3277 493
rect -3311 391 -3277 425
rect -3311 323 -3277 357
rect -3177 521 -3143 540
rect -3177 453 -3143 455
rect -3177 417 -3143 419
rect -3177 332 -3143 351
rect -3019 521 -2985 540
rect -3019 453 -2985 455
rect -3019 417 -2985 419
rect -3019 332 -2985 351
rect -2861 521 -2827 540
rect -2861 453 -2827 455
rect -2861 417 -2827 419
rect -2861 332 -2827 351
rect -2703 521 -2669 540
rect -2703 453 -2669 455
rect -2703 417 -2669 419
rect -2703 332 -2669 351
rect -2545 521 -2511 540
rect -2545 453 -2511 455
rect -2545 417 -2511 419
rect -2545 332 -2511 351
rect -2387 521 -2353 540
rect -2387 453 -2353 455
rect -2387 417 -2353 419
rect -2387 332 -2353 351
rect -2229 521 -2195 540
rect -2229 453 -2195 455
rect -2229 417 -2195 419
rect -2229 332 -2195 351
rect -2071 521 -2037 540
rect -2071 453 -2037 455
rect -2071 417 -2037 419
rect -2071 332 -2037 351
rect -1913 521 -1879 540
rect -1913 453 -1879 455
rect -1913 417 -1879 419
rect -1913 332 -1879 351
rect -1755 521 -1721 540
rect -1755 453 -1721 455
rect -1755 417 -1721 419
rect -1755 332 -1721 351
rect -1597 521 -1563 540
rect -1597 453 -1563 455
rect -1597 417 -1563 419
rect -1597 332 -1563 351
rect -1439 521 -1405 540
rect -1439 453 -1405 455
rect -1439 417 -1405 419
rect -1439 332 -1405 351
rect -1281 521 -1247 540
rect -1281 453 -1247 455
rect -1281 417 -1247 419
rect -1281 332 -1247 351
rect -1123 521 -1089 540
rect -1123 453 -1089 455
rect -1123 417 -1089 419
rect -1123 332 -1089 351
rect -965 521 -931 540
rect -965 453 -931 455
rect -965 417 -931 419
rect -965 332 -931 351
rect -807 521 -773 540
rect -807 453 -773 455
rect -807 417 -773 419
rect -807 332 -773 351
rect -649 521 -615 540
rect -649 453 -615 455
rect -649 417 -615 419
rect -649 332 -615 351
rect -491 521 -457 540
rect -491 453 -457 455
rect -491 417 -457 419
rect -491 332 -457 351
rect -333 521 -299 540
rect -333 453 -299 455
rect -333 417 -299 419
rect -333 332 -299 351
rect -175 521 -141 540
rect -175 453 -141 455
rect -175 417 -141 419
rect -175 332 -141 351
rect -17 521 17 540
rect -17 453 17 455
rect -17 417 17 419
rect -17 332 17 351
rect 141 521 175 540
rect 141 453 175 455
rect 141 417 175 419
rect 141 332 175 351
rect 299 521 333 540
rect 299 453 333 455
rect 299 417 333 419
rect 299 332 333 351
rect 457 521 491 540
rect 457 453 491 455
rect 457 417 491 419
rect 457 332 491 351
rect 615 521 649 540
rect 615 453 649 455
rect 615 417 649 419
rect 615 332 649 351
rect 773 521 807 540
rect 773 453 807 455
rect 773 417 807 419
rect 773 332 807 351
rect 931 521 965 540
rect 931 453 965 455
rect 931 417 965 419
rect 931 332 965 351
rect 1089 521 1123 540
rect 1089 453 1123 455
rect 1089 417 1123 419
rect 1089 332 1123 351
rect 1247 521 1281 540
rect 1247 453 1281 455
rect 1247 417 1281 419
rect 1247 332 1281 351
rect 1405 521 1439 540
rect 1405 453 1439 455
rect 1405 417 1439 419
rect 1405 332 1439 351
rect 1563 521 1597 540
rect 1563 453 1597 455
rect 1563 417 1597 419
rect 1563 332 1597 351
rect 1721 521 1755 540
rect 1721 453 1755 455
rect 1721 417 1755 419
rect 1721 332 1755 351
rect 1879 521 1913 540
rect 1879 453 1913 455
rect 1879 417 1913 419
rect 1879 332 1913 351
rect 2037 521 2071 540
rect 2037 453 2071 455
rect 2037 417 2071 419
rect 2037 332 2071 351
rect 2195 521 2229 540
rect 2195 453 2229 455
rect 2195 417 2229 419
rect 2195 332 2229 351
rect 2353 521 2387 540
rect 2353 453 2387 455
rect 2353 417 2387 419
rect 2353 332 2387 351
rect 2511 521 2545 540
rect 2511 453 2545 455
rect 2511 417 2545 419
rect 2511 332 2545 351
rect 2669 521 2703 540
rect 2669 453 2703 455
rect 2669 417 2703 419
rect 2669 332 2703 351
rect 2827 521 2861 540
rect 2827 453 2861 455
rect 2827 417 2861 419
rect 2827 332 2861 351
rect 2985 521 3019 540
rect 2985 453 3019 455
rect 2985 417 3019 419
rect 2985 332 3019 351
rect 3143 521 3177 540
rect 3143 453 3177 455
rect 3143 417 3177 419
rect 3143 332 3177 351
rect 3277 527 3311 561
rect 3277 459 3311 493
rect 3277 391 3311 425
rect 3277 323 3311 357
rect -3311 255 -3277 289
rect -3131 255 -3098 289
rect -3064 255 -3031 289
rect -2973 255 -2940 289
rect -2906 255 -2873 289
rect -2815 255 -2782 289
rect -2748 255 -2715 289
rect -2657 255 -2624 289
rect -2590 255 -2557 289
rect -2499 255 -2466 289
rect -2432 255 -2399 289
rect -2341 255 -2308 289
rect -2274 255 -2241 289
rect -2183 255 -2150 289
rect -2116 255 -2083 289
rect -2025 255 -1992 289
rect -1958 255 -1925 289
rect -1867 255 -1834 289
rect -1800 255 -1767 289
rect -1709 255 -1676 289
rect -1642 255 -1609 289
rect -1551 255 -1518 289
rect -1484 255 -1451 289
rect -1393 255 -1360 289
rect -1326 255 -1293 289
rect -1235 255 -1202 289
rect -1168 255 -1135 289
rect -1077 255 -1044 289
rect -1010 255 -977 289
rect -919 255 -886 289
rect -852 255 -819 289
rect -761 255 -728 289
rect -694 255 -661 289
rect -603 255 -570 289
rect -536 255 -503 289
rect -445 255 -412 289
rect -378 255 -345 289
rect -287 255 -254 289
rect -220 255 -187 289
rect -129 255 -96 289
rect -62 255 -29 289
rect 29 255 62 289
rect 96 255 129 289
rect 187 255 220 289
rect 254 255 287 289
rect 345 255 378 289
rect 412 255 445 289
rect 503 255 536 289
rect 570 255 603 289
rect 661 255 694 289
rect 728 255 761 289
rect 819 255 852 289
rect 886 255 919 289
rect 977 255 1010 289
rect 1044 255 1077 289
rect 1135 255 1168 289
rect 1202 255 1235 289
rect 1293 255 1326 289
rect 1360 255 1393 289
rect 1451 255 1484 289
rect 1518 255 1551 289
rect 1609 255 1642 289
rect 1676 255 1709 289
rect 1767 255 1800 289
rect 1834 255 1867 289
rect 1925 255 1958 289
rect 1992 255 2025 289
rect 2083 255 2116 289
rect 2150 255 2183 289
rect 2241 255 2274 289
rect 2308 255 2341 289
rect 2399 255 2432 289
rect 2466 255 2499 289
rect 2557 255 2590 289
rect 2624 255 2657 289
rect 2715 255 2748 289
rect 2782 255 2815 289
rect 2873 255 2906 289
rect 2940 255 2973 289
rect 3031 255 3064 289
rect 3098 255 3131 289
rect 3277 255 3311 289
rect -3311 187 -3277 221
rect 3277 187 3311 221
rect -3311 119 -3277 153
rect -3131 147 -3098 181
rect -3064 147 -3031 181
rect -2973 147 -2940 181
rect -2906 147 -2873 181
rect -2815 147 -2782 181
rect -2748 147 -2715 181
rect -2657 147 -2624 181
rect -2590 147 -2557 181
rect -2499 147 -2466 181
rect -2432 147 -2399 181
rect -2341 147 -2308 181
rect -2274 147 -2241 181
rect -2183 147 -2150 181
rect -2116 147 -2083 181
rect -2025 147 -1992 181
rect -1958 147 -1925 181
rect -1867 147 -1834 181
rect -1800 147 -1767 181
rect -1709 147 -1676 181
rect -1642 147 -1609 181
rect -1551 147 -1518 181
rect -1484 147 -1451 181
rect -1393 147 -1360 181
rect -1326 147 -1293 181
rect -1235 147 -1202 181
rect -1168 147 -1135 181
rect -1077 147 -1044 181
rect -1010 147 -977 181
rect -919 147 -886 181
rect -852 147 -819 181
rect -761 147 -728 181
rect -694 147 -661 181
rect -603 147 -570 181
rect -536 147 -503 181
rect -445 147 -412 181
rect -378 147 -345 181
rect -287 147 -254 181
rect -220 147 -187 181
rect -129 147 -96 181
rect -62 147 -29 181
rect 29 147 62 181
rect 96 147 129 181
rect 187 147 220 181
rect 254 147 287 181
rect 345 147 378 181
rect 412 147 445 181
rect 503 147 536 181
rect 570 147 603 181
rect 661 147 694 181
rect 728 147 761 181
rect 819 147 852 181
rect 886 147 919 181
rect 977 147 1010 181
rect 1044 147 1077 181
rect 1135 147 1168 181
rect 1202 147 1235 181
rect 1293 147 1326 181
rect 1360 147 1393 181
rect 1451 147 1484 181
rect 1518 147 1551 181
rect 1609 147 1642 181
rect 1676 147 1709 181
rect 1767 147 1800 181
rect 1834 147 1867 181
rect 1925 147 1958 181
rect 1992 147 2025 181
rect 2083 147 2116 181
rect 2150 147 2183 181
rect 2241 147 2274 181
rect 2308 147 2341 181
rect 2399 147 2432 181
rect 2466 147 2499 181
rect 2557 147 2590 181
rect 2624 147 2657 181
rect 2715 147 2748 181
rect 2782 147 2815 181
rect 2873 147 2906 181
rect 2940 147 2973 181
rect 3031 147 3064 181
rect 3098 147 3131 181
rect 3277 119 3311 153
rect -3311 51 -3277 85
rect -3311 -17 -3277 17
rect -3311 -85 -3277 -51
rect -3177 85 -3143 104
rect -3177 17 -3143 19
rect -3177 -19 -3143 -17
rect -3177 -104 -3143 -85
rect -3019 85 -2985 104
rect -3019 17 -2985 19
rect -3019 -19 -2985 -17
rect -3019 -104 -2985 -85
rect -2861 85 -2827 104
rect -2861 17 -2827 19
rect -2861 -19 -2827 -17
rect -2861 -104 -2827 -85
rect -2703 85 -2669 104
rect -2703 17 -2669 19
rect -2703 -19 -2669 -17
rect -2703 -104 -2669 -85
rect -2545 85 -2511 104
rect -2545 17 -2511 19
rect -2545 -19 -2511 -17
rect -2545 -104 -2511 -85
rect -2387 85 -2353 104
rect -2387 17 -2353 19
rect -2387 -19 -2353 -17
rect -2387 -104 -2353 -85
rect -2229 85 -2195 104
rect -2229 17 -2195 19
rect -2229 -19 -2195 -17
rect -2229 -104 -2195 -85
rect -2071 85 -2037 104
rect -2071 17 -2037 19
rect -2071 -19 -2037 -17
rect -2071 -104 -2037 -85
rect -1913 85 -1879 104
rect -1913 17 -1879 19
rect -1913 -19 -1879 -17
rect -1913 -104 -1879 -85
rect -1755 85 -1721 104
rect -1755 17 -1721 19
rect -1755 -19 -1721 -17
rect -1755 -104 -1721 -85
rect -1597 85 -1563 104
rect -1597 17 -1563 19
rect -1597 -19 -1563 -17
rect -1597 -104 -1563 -85
rect -1439 85 -1405 104
rect -1439 17 -1405 19
rect -1439 -19 -1405 -17
rect -1439 -104 -1405 -85
rect -1281 85 -1247 104
rect -1281 17 -1247 19
rect -1281 -19 -1247 -17
rect -1281 -104 -1247 -85
rect -1123 85 -1089 104
rect -1123 17 -1089 19
rect -1123 -19 -1089 -17
rect -1123 -104 -1089 -85
rect -965 85 -931 104
rect -965 17 -931 19
rect -965 -19 -931 -17
rect -965 -104 -931 -85
rect -807 85 -773 104
rect -807 17 -773 19
rect -807 -19 -773 -17
rect -807 -104 -773 -85
rect -649 85 -615 104
rect -649 17 -615 19
rect -649 -19 -615 -17
rect -649 -104 -615 -85
rect -491 85 -457 104
rect -491 17 -457 19
rect -491 -19 -457 -17
rect -491 -104 -457 -85
rect -333 85 -299 104
rect -333 17 -299 19
rect -333 -19 -299 -17
rect -333 -104 -299 -85
rect -175 85 -141 104
rect -175 17 -141 19
rect -175 -19 -141 -17
rect -175 -104 -141 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 141 85 175 104
rect 141 17 175 19
rect 141 -19 175 -17
rect 141 -104 175 -85
rect 299 85 333 104
rect 299 17 333 19
rect 299 -19 333 -17
rect 299 -104 333 -85
rect 457 85 491 104
rect 457 17 491 19
rect 457 -19 491 -17
rect 457 -104 491 -85
rect 615 85 649 104
rect 615 17 649 19
rect 615 -19 649 -17
rect 615 -104 649 -85
rect 773 85 807 104
rect 773 17 807 19
rect 773 -19 807 -17
rect 773 -104 807 -85
rect 931 85 965 104
rect 931 17 965 19
rect 931 -19 965 -17
rect 931 -104 965 -85
rect 1089 85 1123 104
rect 1089 17 1123 19
rect 1089 -19 1123 -17
rect 1089 -104 1123 -85
rect 1247 85 1281 104
rect 1247 17 1281 19
rect 1247 -19 1281 -17
rect 1247 -104 1281 -85
rect 1405 85 1439 104
rect 1405 17 1439 19
rect 1405 -19 1439 -17
rect 1405 -104 1439 -85
rect 1563 85 1597 104
rect 1563 17 1597 19
rect 1563 -19 1597 -17
rect 1563 -104 1597 -85
rect 1721 85 1755 104
rect 1721 17 1755 19
rect 1721 -19 1755 -17
rect 1721 -104 1755 -85
rect 1879 85 1913 104
rect 1879 17 1913 19
rect 1879 -19 1913 -17
rect 1879 -104 1913 -85
rect 2037 85 2071 104
rect 2037 17 2071 19
rect 2037 -19 2071 -17
rect 2037 -104 2071 -85
rect 2195 85 2229 104
rect 2195 17 2229 19
rect 2195 -19 2229 -17
rect 2195 -104 2229 -85
rect 2353 85 2387 104
rect 2353 17 2387 19
rect 2353 -19 2387 -17
rect 2353 -104 2387 -85
rect 2511 85 2545 104
rect 2511 17 2545 19
rect 2511 -19 2545 -17
rect 2511 -104 2545 -85
rect 2669 85 2703 104
rect 2669 17 2703 19
rect 2669 -19 2703 -17
rect 2669 -104 2703 -85
rect 2827 85 2861 104
rect 2827 17 2861 19
rect 2827 -19 2861 -17
rect 2827 -104 2861 -85
rect 2985 85 3019 104
rect 2985 17 3019 19
rect 2985 -19 3019 -17
rect 2985 -104 3019 -85
rect 3143 85 3177 104
rect 3143 17 3177 19
rect 3143 -19 3177 -17
rect 3143 -104 3177 -85
rect 3277 51 3311 85
rect 3277 -17 3311 17
rect 3277 -85 3311 -51
rect -3311 -153 -3277 -119
rect -3131 -181 -3098 -147
rect -3064 -181 -3031 -147
rect -2973 -181 -2940 -147
rect -2906 -181 -2873 -147
rect -2815 -181 -2782 -147
rect -2748 -181 -2715 -147
rect -2657 -181 -2624 -147
rect -2590 -181 -2557 -147
rect -2499 -181 -2466 -147
rect -2432 -181 -2399 -147
rect -2341 -181 -2308 -147
rect -2274 -181 -2241 -147
rect -2183 -181 -2150 -147
rect -2116 -181 -2083 -147
rect -2025 -181 -1992 -147
rect -1958 -181 -1925 -147
rect -1867 -181 -1834 -147
rect -1800 -181 -1767 -147
rect -1709 -181 -1676 -147
rect -1642 -181 -1609 -147
rect -1551 -181 -1518 -147
rect -1484 -181 -1451 -147
rect -1393 -181 -1360 -147
rect -1326 -181 -1293 -147
rect -1235 -181 -1202 -147
rect -1168 -181 -1135 -147
rect -1077 -181 -1044 -147
rect -1010 -181 -977 -147
rect -919 -181 -886 -147
rect -852 -181 -819 -147
rect -761 -181 -728 -147
rect -694 -181 -661 -147
rect -603 -181 -570 -147
rect -536 -181 -503 -147
rect -445 -181 -412 -147
rect -378 -181 -345 -147
rect -287 -181 -254 -147
rect -220 -181 -187 -147
rect -129 -181 -96 -147
rect -62 -181 -29 -147
rect 29 -181 62 -147
rect 96 -181 129 -147
rect 187 -181 220 -147
rect 254 -181 287 -147
rect 345 -181 378 -147
rect 412 -181 445 -147
rect 503 -181 536 -147
rect 570 -181 603 -147
rect 661 -181 694 -147
rect 728 -181 761 -147
rect 819 -181 852 -147
rect 886 -181 919 -147
rect 977 -181 1010 -147
rect 1044 -181 1077 -147
rect 1135 -181 1168 -147
rect 1202 -181 1235 -147
rect 1293 -181 1326 -147
rect 1360 -181 1393 -147
rect 1451 -181 1484 -147
rect 1518 -181 1551 -147
rect 1609 -181 1642 -147
rect 1676 -181 1709 -147
rect 1767 -181 1800 -147
rect 1834 -181 1867 -147
rect 1925 -181 1958 -147
rect 1992 -181 2025 -147
rect 2083 -181 2116 -147
rect 2150 -181 2183 -147
rect 2241 -181 2274 -147
rect 2308 -181 2341 -147
rect 2399 -181 2432 -147
rect 2466 -181 2499 -147
rect 2557 -181 2590 -147
rect 2624 -181 2657 -147
rect 2715 -181 2748 -147
rect 2782 -181 2815 -147
rect 2873 -181 2906 -147
rect 2940 -181 2973 -147
rect 3031 -181 3064 -147
rect 3098 -181 3131 -147
rect 3277 -153 3311 -119
rect -3311 -221 -3277 -187
rect 3277 -221 3311 -187
rect -3311 -289 -3277 -255
rect -3131 -289 -3098 -255
rect -3064 -289 -3031 -255
rect -2973 -289 -2940 -255
rect -2906 -289 -2873 -255
rect -2815 -289 -2782 -255
rect -2748 -289 -2715 -255
rect -2657 -289 -2624 -255
rect -2590 -289 -2557 -255
rect -2499 -289 -2466 -255
rect -2432 -289 -2399 -255
rect -2341 -289 -2308 -255
rect -2274 -289 -2241 -255
rect -2183 -289 -2150 -255
rect -2116 -289 -2083 -255
rect -2025 -289 -1992 -255
rect -1958 -289 -1925 -255
rect -1867 -289 -1834 -255
rect -1800 -289 -1767 -255
rect -1709 -289 -1676 -255
rect -1642 -289 -1609 -255
rect -1551 -289 -1518 -255
rect -1484 -289 -1451 -255
rect -1393 -289 -1360 -255
rect -1326 -289 -1293 -255
rect -1235 -289 -1202 -255
rect -1168 -289 -1135 -255
rect -1077 -289 -1044 -255
rect -1010 -289 -977 -255
rect -919 -289 -886 -255
rect -852 -289 -819 -255
rect -761 -289 -728 -255
rect -694 -289 -661 -255
rect -603 -289 -570 -255
rect -536 -289 -503 -255
rect -445 -289 -412 -255
rect -378 -289 -345 -255
rect -287 -289 -254 -255
rect -220 -289 -187 -255
rect -129 -289 -96 -255
rect -62 -289 -29 -255
rect 29 -289 62 -255
rect 96 -289 129 -255
rect 187 -289 220 -255
rect 254 -289 287 -255
rect 345 -289 378 -255
rect 412 -289 445 -255
rect 503 -289 536 -255
rect 570 -289 603 -255
rect 661 -289 694 -255
rect 728 -289 761 -255
rect 819 -289 852 -255
rect 886 -289 919 -255
rect 977 -289 1010 -255
rect 1044 -289 1077 -255
rect 1135 -289 1168 -255
rect 1202 -289 1235 -255
rect 1293 -289 1326 -255
rect 1360 -289 1393 -255
rect 1451 -289 1484 -255
rect 1518 -289 1551 -255
rect 1609 -289 1642 -255
rect 1676 -289 1709 -255
rect 1767 -289 1800 -255
rect 1834 -289 1867 -255
rect 1925 -289 1958 -255
rect 1992 -289 2025 -255
rect 2083 -289 2116 -255
rect 2150 -289 2183 -255
rect 2241 -289 2274 -255
rect 2308 -289 2341 -255
rect 2399 -289 2432 -255
rect 2466 -289 2499 -255
rect 2557 -289 2590 -255
rect 2624 -289 2657 -255
rect 2715 -289 2748 -255
rect 2782 -289 2815 -255
rect 2873 -289 2906 -255
rect 2940 -289 2973 -255
rect 3031 -289 3064 -255
rect 3098 -289 3131 -255
rect 3277 -289 3311 -255
rect -3311 -357 -3277 -323
rect -3311 -425 -3277 -391
rect -3311 -493 -3277 -459
rect -3311 -561 -3277 -527
rect -3177 -351 -3143 -332
rect -3177 -419 -3143 -417
rect -3177 -455 -3143 -453
rect -3177 -540 -3143 -521
rect -3019 -351 -2985 -332
rect -3019 -419 -2985 -417
rect -3019 -455 -2985 -453
rect -3019 -540 -2985 -521
rect -2861 -351 -2827 -332
rect -2861 -419 -2827 -417
rect -2861 -455 -2827 -453
rect -2861 -540 -2827 -521
rect -2703 -351 -2669 -332
rect -2703 -419 -2669 -417
rect -2703 -455 -2669 -453
rect -2703 -540 -2669 -521
rect -2545 -351 -2511 -332
rect -2545 -419 -2511 -417
rect -2545 -455 -2511 -453
rect -2545 -540 -2511 -521
rect -2387 -351 -2353 -332
rect -2387 -419 -2353 -417
rect -2387 -455 -2353 -453
rect -2387 -540 -2353 -521
rect -2229 -351 -2195 -332
rect -2229 -419 -2195 -417
rect -2229 -455 -2195 -453
rect -2229 -540 -2195 -521
rect -2071 -351 -2037 -332
rect -2071 -419 -2037 -417
rect -2071 -455 -2037 -453
rect -2071 -540 -2037 -521
rect -1913 -351 -1879 -332
rect -1913 -419 -1879 -417
rect -1913 -455 -1879 -453
rect -1913 -540 -1879 -521
rect -1755 -351 -1721 -332
rect -1755 -419 -1721 -417
rect -1755 -455 -1721 -453
rect -1755 -540 -1721 -521
rect -1597 -351 -1563 -332
rect -1597 -419 -1563 -417
rect -1597 -455 -1563 -453
rect -1597 -540 -1563 -521
rect -1439 -351 -1405 -332
rect -1439 -419 -1405 -417
rect -1439 -455 -1405 -453
rect -1439 -540 -1405 -521
rect -1281 -351 -1247 -332
rect -1281 -419 -1247 -417
rect -1281 -455 -1247 -453
rect -1281 -540 -1247 -521
rect -1123 -351 -1089 -332
rect -1123 -419 -1089 -417
rect -1123 -455 -1089 -453
rect -1123 -540 -1089 -521
rect -965 -351 -931 -332
rect -965 -419 -931 -417
rect -965 -455 -931 -453
rect -965 -540 -931 -521
rect -807 -351 -773 -332
rect -807 -419 -773 -417
rect -807 -455 -773 -453
rect -807 -540 -773 -521
rect -649 -351 -615 -332
rect -649 -419 -615 -417
rect -649 -455 -615 -453
rect -649 -540 -615 -521
rect -491 -351 -457 -332
rect -491 -419 -457 -417
rect -491 -455 -457 -453
rect -491 -540 -457 -521
rect -333 -351 -299 -332
rect -333 -419 -299 -417
rect -333 -455 -299 -453
rect -333 -540 -299 -521
rect -175 -351 -141 -332
rect -175 -419 -141 -417
rect -175 -455 -141 -453
rect -175 -540 -141 -521
rect -17 -351 17 -332
rect -17 -419 17 -417
rect -17 -455 17 -453
rect -17 -540 17 -521
rect 141 -351 175 -332
rect 141 -419 175 -417
rect 141 -455 175 -453
rect 141 -540 175 -521
rect 299 -351 333 -332
rect 299 -419 333 -417
rect 299 -455 333 -453
rect 299 -540 333 -521
rect 457 -351 491 -332
rect 457 -419 491 -417
rect 457 -455 491 -453
rect 457 -540 491 -521
rect 615 -351 649 -332
rect 615 -419 649 -417
rect 615 -455 649 -453
rect 615 -540 649 -521
rect 773 -351 807 -332
rect 773 -419 807 -417
rect 773 -455 807 -453
rect 773 -540 807 -521
rect 931 -351 965 -332
rect 931 -419 965 -417
rect 931 -455 965 -453
rect 931 -540 965 -521
rect 1089 -351 1123 -332
rect 1089 -419 1123 -417
rect 1089 -455 1123 -453
rect 1089 -540 1123 -521
rect 1247 -351 1281 -332
rect 1247 -419 1281 -417
rect 1247 -455 1281 -453
rect 1247 -540 1281 -521
rect 1405 -351 1439 -332
rect 1405 -419 1439 -417
rect 1405 -455 1439 -453
rect 1405 -540 1439 -521
rect 1563 -351 1597 -332
rect 1563 -419 1597 -417
rect 1563 -455 1597 -453
rect 1563 -540 1597 -521
rect 1721 -351 1755 -332
rect 1721 -419 1755 -417
rect 1721 -455 1755 -453
rect 1721 -540 1755 -521
rect 1879 -351 1913 -332
rect 1879 -419 1913 -417
rect 1879 -455 1913 -453
rect 1879 -540 1913 -521
rect 2037 -351 2071 -332
rect 2037 -419 2071 -417
rect 2037 -455 2071 -453
rect 2037 -540 2071 -521
rect 2195 -351 2229 -332
rect 2195 -419 2229 -417
rect 2195 -455 2229 -453
rect 2195 -540 2229 -521
rect 2353 -351 2387 -332
rect 2353 -419 2387 -417
rect 2353 -455 2387 -453
rect 2353 -540 2387 -521
rect 2511 -351 2545 -332
rect 2511 -419 2545 -417
rect 2511 -455 2545 -453
rect 2511 -540 2545 -521
rect 2669 -351 2703 -332
rect 2669 -419 2703 -417
rect 2669 -455 2703 -453
rect 2669 -540 2703 -521
rect 2827 -351 2861 -332
rect 2827 -419 2861 -417
rect 2827 -455 2861 -453
rect 2827 -540 2861 -521
rect 2985 -351 3019 -332
rect 2985 -419 3019 -417
rect 2985 -455 3019 -453
rect 2985 -540 3019 -521
rect 3143 -351 3177 -332
rect 3143 -419 3177 -417
rect 3143 -455 3177 -453
rect 3143 -540 3177 -521
rect 3277 -357 3311 -323
rect 3277 -425 3311 -391
rect 3277 -493 3311 -459
rect 3277 -561 3311 -527
rect -3311 -629 -3277 -595
rect -3131 -617 -3098 -583
rect -3064 -617 -3031 -583
rect -2973 -617 -2940 -583
rect -2906 -617 -2873 -583
rect -2815 -617 -2782 -583
rect -2748 -617 -2715 -583
rect -2657 -617 -2624 -583
rect -2590 -617 -2557 -583
rect -2499 -617 -2466 -583
rect -2432 -617 -2399 -583
rect -2341 -617 -2308 -583
rect -2274 -617 -2241 -583
rect -2183 -617 -2150 -583
rect -2116 -617 -2083 -583
rect -2025 -617 -1992 -583
rect -1958 -617 -1925 -583
rect -1867 -617 -1834 -583
rect -1800 -617 -1767 -583
rect -1709 -617 -1676 -583
rect -1642 -617 -1609 -583
rect -1551 -617 -1518 -583
rect -1484 -617 -1451 -583
rect -1393 -617 -1360 -583
rect -1326 -617 -1293 -583
rect -1235 -617 -1202 -583
rect -1168 -617 -1135 -583
rect -1077 -617 -1044 -583
rect -1010 -617 -977 -583
rect -919 -617 -886 -583
rect -852 -617 -819 -583
rect -761 -617 -728 -583
rect -694 -617 -661 -583
rect -603 -617 -570 -583
rect -536 -617 -503 -583
rect -445 -617 -412 -583
rect -378 -617 -345 -583
rect -287 -617 -254 -583
rect -220 -617 -187 -583
rect -129 -617 -96 -583
rect -62 -617 -29 -583
rect 29 -617 62 -583
rect 96 -617 129 -583
rect 187 -617 220 -583
rect 254 -617 287 -583
rect 345 -617 378 -583
rect 412 -617 445 -583
rect 503 -617 536 -583
rect 570 -617 603 -583
rect 661 -617 694 -583
rect 728 -617 761 -583
rect 819 -617 852 -583
rect 886 -617 919 -583
rect 977 -617 1010 -583
rect 1044 -617 1077 -583
rect 1135 -617 1168 -583
rect 1202 -617 1235 -583
rect 1293 -617 1326 -583
rect 1360 -617 1393 -583
rect 1451 -617 1484 -583
rect 1518 -617 1551 -583
rect 1609 -617 1642 -583
rect 1676 -617 1709 -583
rect 1767 -617 1800 -583
rect 1834 -617 1867 -583
rect 1925 -617 1958 -583
rect 1992 -617 2025 -583
rect 2083 -617 2116 -583
rect 2150 -617 2183 -583
rect 2241 -617 2274 -583
rect 2308 -617 2341 -583
rect 2399 -617 2432 -583
rect 2466 -617 2499 -583
rect 2557 -617 2590 -583
rect 2624 -617 2657 -583
rect 2715 -617 2748 -583
rect 2782 -617 2815 -583
rect 2873 -617 2906 -583
rect 2940 -617 2973 -583
rect 3031 -617 3064 -583
rect 3098 -617 3131 -583
rect -3311 -697 -3277 -663
rect 3277 -629 3311 -595
rect -3131 -725 -3098 -691
rect -3064 -725 -3031 -691
rect -2973 -725 -2940 -691
rect -2906 -725 -2873 -691
rect -2815 -725 -2782 -691
rect -2748 -725 -2715 -691
rect -2657 -725 -2624 -691
rect -2590 -725 -2557 -691
rect -2499 -725 -2466 -691
rect -2432 -725 -2399 -691
rect -2341 -725 -2308 -691
rect -2274 -725 -2241 -691
rect -2183 -725 -2150 -691
rect -2116 -725 -2083 -691
rect -2025 -725 -1992 -691
rect -1958 -725 -1925 -691
rect -1867 -725 -1834 -691
rect -1800 -725 -1767 -691
rect -1709 -725 -1676 -691
rect -1642 -725 -1609 -691
rect -1551 -725 -1518 -691
rect -1484 -725 -1451 -691
rect -1393 -725 -1360 -691
rect -1326 -725 -1293 -691
rect -1235 -725 -1202 -691
rect -1168 -725 -1135 -691
rect -1077 -725 -1044 -691
rect -1010 -725 -977 -691
rect -919 -725 -886 -691
rect -852 -725 -819 -691
rect -761 -725 -728 -691
rect -694 -725 -661 -691
rect -603 -725 -570 -691
rect -536 -725 -503 -691
rect -445 -725 -412 -691
rect -378 -725 -345 -691
rect -287 -725 -254 -691
rect -220 -725 -187 -691
rect -129 -725 -96 -691
rect -62 -725 -29 -691
rect 29 -725 62 -691
rect 96 -725 129 -691
rect 187 -725 220 -691
rect 254 -725 287 -691
rect 345 -725 378 -691
rect 412 -725 445 -691
rect 503 -725 536 -691
rect 570 -725 603 -691
rect 661 -725 694 -691
rect 728 -725 761 -691
rect 819 -725 852 -691
rect 886 -725 919 -691
rect 977 -725 1010 -691
rect 1044 -725 1077 -691
rect 1135 -725 1168 -691
rect 1202 -725 1235 -691
rect 1293 -725 1326 -691
rect 1360 -725 1393 -691
rect 1451 -725 1484 -691
rect 1518 -725 1551 -691
rect 1609 -725 1642 -691
rect 1676 -725 1709 -691
rect 1767 -725 1800 -691
rect 1834 -725 1867 -691
rect 1925 -725 1958 -691
rect 1992 -725 2025 -691
rect 2083 -725 2116 -691
rect 2150 -725 2183 -691
rect 2241 -725 2274 -691
rect 2308 -725 2341 -691
rect 2399 -725 2432 -691
rect 2466 -725 2499 -691
rect 2557 -725 2590 -691
rect 2624 -725 2657 -691
rect 2715 -725 2748 -691
rect 2782 -725 2815 -691
rect 2873 -725 2906 -691
rect 2940 -725 2973 -691
rect 3031 -725 3064 -691
rect 3098 -725 3131 -691
rect 3277 -697 3311 -663
rect -3311 -765 -3277 -731
rect 3277 -765 3311 -731
rect -3311 -833 -3277 -799
rect -3311 -901 -3277 -867
rect -3311 -969 -3277 -935
rect -3177 -787 -3143 -768
rect -3177 -855 -3143 -853
rect -3177 -891 -3143 -889
rect -3177 -976 -3143 -957
rect -3019 -787 -2985 -768
rect -3019 -855 -2985 -853
rect -3019 -891 -2985 -889
rect -3019 -976 -2985 -957
rect -2861 -787 -2827 -768
rect -2861 -855 -2827 -853
rect -2861 -891 -2827 -889
rect -2861 -976 -2827 -957
rect -2703 -787 -2669 -768
rect -2703 -855 -2669 -853
rect -2703 -891 -2669 -889
rect -2703 -976 -2669 -957
rect -2545 -787 -2511 -768
rect -2545 -855 -2511 -853
rect -2545 -891 -2511 -889
rect -2545 -976 -2511 -957
rect -2387 -787 -2353 -768
rect -2387 -855 -2353 -853
rect -2387 -891 -2353 -889
rect -2387 -976 -2353 -957
rect -2229 -787 -2195 -768
rect -2229 -855 -2195 -853
rect -2229 -891 -2195 -889
rect -2229 -976 -2195 -957
rect -2071 -787 -2037 -768
rect -2071 -855 -2037 -853
rect -2071 -891 -2037 -889
rect -2071 -976 -2037 -957
rect -1913 -787 -1879 -768
rect -1913 -855 -1879 -853
rect -1913 -891 -1879 -889
rect -1913 -976 -1879 -957
rect -1755 -787 -1721 -768
rect -1755 -855 -1721 -853
rect -1755 -891 -1721 -889
rect -1755 -976 -1721 -957
rect -1597 -787 -1563 -768
rect -1597 -855 -1563 -853
rect -1597 -891 -1563 -889
rect -1597 -976 -1563 -957
rect -1439 -787 -1405 -768
rect -1439 -855 -1405 -853
rect -1439 -891 -1405 -889
rect -1439 -976 -1405 -957
rect -1281 -787 -1247 -768
rect -1281 -855 -1247 -853
rect -1281 -891 -1247 -889
rect -1281 -976 -1247 -957
rect -1123 -787 -1089 -768
rect -1123 -855 -1089 -853
rect -1123 -891 -1089 -889
rect -1123 -976 -1089 -957
rect -965 -787 -931 -768
rect -965 -855 -931 -853
rect -965 -891 -931 -889
rect -965 -976 -931 -957
rect -807 -787 -773 -768
rect -807 -855 -773 -853
rect -807 -891 -773 -889
rect -807 -976 -773 -957
rect -649 -787 -615 -768
rect -649 -855 -615 -853
rect -649 -891 -615 -889
rect -649 -976 -615 -957
rect -491 -787 -457 -768
rect -491 -855 -457 -853
rect -491 -891 -457 -889
rect -491 -976 -457 -957
rect -333 -787 -299 -768
rect -333 -855 -299 -853
rect -333 -891 -299 -889
rect -333 -976 -299 -957
rect -175 -787 -141 -768
rect -175 -855 -141 -853
rect -175 -891 -141 -889
rect -175 -976 -141 -957
rect -17 -787 17 -768
rect -17 -855 17 -853
rect -17 -891 17 -889
rect -17 -976 17 -957
rect 141 -787 175 -768
rect 141 -855 175 -853
rect 141 -891 175 -889
rect 141 -976 175 -957
rect 299 -787 333 -768
rect 299 -855 333 -853
rect 299 -891 333 -889
rect 299 -976 333 -957
rect 457 -787 491 -768
rect 457 -855 491 -853
rect 457 -891 491 -889
rect 457 -976 491 -957
rect 615 -787 649 -768
rect 615 -855 649 -853
rect 615 -891 649 -889
rect 615 -976 649 -957
rect 773 -787 807 -768
rect 773 -855 807 -853
rect 773 -891 807 -889
rect 773 -976 807 -957
rect 931 -787 965 -768
rect 931 -855 965 -853
rect 931 -891 965 -889
rect 931 -976 965 -957
rect 1089 -787 1123 -768
rect 1089 -855 1123 -853
rect 1089 -891 1123 -889
rect 1089 -976 1123 -957
rect 1247 -787 1281 -768
rect 1247 -855 1281 -853
rect 1247 -891 1281 -889
rect 1247 -976 1281 -957
rect 1405 -787 1439 -768
rect 1405 -855 1439 -853
rect 1405 -891 1439 -889
rect 1405 -976 1439 -957
rect 1563 -787 1597 -768
rect 1563 -855 1597 -853
rect 1563 -891 1597 -889
rect 1563 -976 1597 -957
rect 1721 -787 1755 -768
rect 1721 -855 1755 -853
rect 1721 -891 1755 -889
rect 1721 -976 1755 -957
rect 1879 -787 1913 -768
rect 1879 -855 1913 -853
rect 1879 -891 1913 -889
rect 1879 -976 1913 -957
rect 2037 -787 2071 -768
rect 2037 -855 2071 -853
rect 2037 -891 2071 -889
rect 2037 -976 2071 -957
rect 2195 -787 2229 -768
rect 2195 -855 2229 -853
rect 2195 -891 2229 -889
rect 2195 -976 2229 -957
rect 2353 -787 2387 -768
rect 2353 -855 2387 -853
rect 2353 -891 2387 -889
rect 2353 -976 2387 -957
rect 2511 -787 2545 -768
rect 2511 -855 2545 -853
rect 2511 -891 2545 -889
rect 2511 -976 2545 -957
rect 2669 -787 2703 -768
rect 2669 -855 2703 -853
rect 2669 -891 2703 -889
rect 2669 -976 2703 -957
rect 2827 -787 2861 -768
rect 2827 -855 2861 -853
rect 2827 -891 2861 -889
rect 2827 -976 2861 -957
rect 2985 -787 3019 -768
rect 2985 -855 3019 -853
rect 2985 -891 3019 -889
rect 2985 -976 3019 -957
rect 3143 -787 3177 -768
rect 3143 -855 3177 -853
rect 3143 -891 3177 -889
rect 3143 -976 3177 -957
rect 3277 -833 3311 -799
rect 3277 -901 3311 -867
rect 3277 -969 3311 -935
rect -3311 -1037 -3277 -1003
rect -3131 -1053 -3098 -1019
rect -3064 -1053 -3031 -1019
rect -2973 -1053 -2940 -1019
rect -2906 -1053 -2873 -1019
rect -2815 -1053 -2782 -1019
rect -2748 -1053 -2715 -1019
rect -2657 -1053 -2624 -1019
rect -2590 -1053 -2557 -1019
rect -2499 -1053 -2466 -1019
rect -2432 -1053 -2399 -1019
rect -2341 -1053 -2308 -1019
rect -2274 -1053 -2241 -1019
rect -2183 -1053 -2150 -1019
rect -2116 -1053 -2083 -1019
rect -2025 -1053 -1992 -1019
rect -1958 -1053 -1925 -1019
rect -1867 -1053 -1834 -1019
rect -1800 -1053 -1767 -1019
rect -1709 -1053 -1676 -1019
rect -1642 -1053 -1609 -1019
rect -1551 -1053 -1518 -1019
rect -1484 -1053 -1451 -1019
rect -1393 -1053 -1360 -1019
rect -1326 -1053 -1293 -1019
rect -1235 -1053 -1202 -1019
rect -1168 -1053 -1135 -1019
rect -1077 -1053 -1044 -1019
rect -1010 -1053 -977 -1019
rect -919 -1053 -886 -1019
rect -852 -1053 -819 -1019
rect -761 -1053 -728 -1019
rect -694 -1053 -661 -1019
rect -603 -1053 -570 -1019
rect -536 -1053 -503 -1019
rect -445 -1053 -412 -1019
rect -378 -1053 -345 -1019
rect -287 -1053 -254 -1019
rect -220 -1053 -187 -1019
rect -129 -1053 -96 -1019
rect -62 -1053 -29 -1019
rect 29 -1053 62 -1019
rect 96 -1053 129 -1019
rect 187 -1053 220 -1019
rect 254 -1053 287 -1019
rect 345 -1053 378 -1019
rect 412 -1053 445 -1019
rect 503 -1053 536 -1019
rect 570 -1053 603 -1019
rect 661 -1053 694 -1019
rect 728 -1053 761 -1019
rect 819 -1053 852 -1019
rect 886 -1053 919 -1019
rect 977 -1053 1010 -1019
rect 1044 -1053 1077 -1019
rect 1135 -1053 1168 -1019
rect 1202 -1053 1235 -1019
rect 1293 -1053 1326 -1019
rect 1360 -1053 1393 -1019
rect 1451 -1053 1484 -1019
rect 1518 -1053 1551 -1019
rect 1609 -1053 1642 -1019
rect 1676 -1053 1709 -1019
rect 1767 -1053 1800 -1019
rect 1834 -1053 1867 -1019
rect 1925 -1053 1958 -1019
rect 1992 -1053 2025 -1019
rect 2083 -1053 2116 -1019
rect 2150 -1053 2183 -1019
rect 2241 -1053 2274 -1019
rect 2308 -1053 2341 -1019
rect 2399 -1053 2432 -1019
rect 2466 -1053 2499 -1019
rect 2557 -1053 2590 -1019
rect 2624 -1053 2657 -1019
rect 2715 -1053 2748 -1019
rect 2782 -1053 2815 -1019
rect 2873 -1053 2906 -1019
rect 2940 -1053 2973 -1019
rect 3031 -1053 3064 -1019
rect 3098 -1053 3131 -1019
rect 3277 -1037 3311 -1003
rect -3311 -1157 -3277 -1071
rect 3277 -1157 3311 -1071
rect -3311 -1191 -3213 -1157
rect -3179 -1191 -3145 -1157
rect -3111 -1191 -3077 -1157
rect -3043 -1191 -3009 -1157
rect -2975 -1191 -2941 -1157
rect -2907 -1191 -2873 -1157
rect -2839 -1191 -2805 -1157
rect -2771 -1191 -2737 -1157
rect -2703 -1191 -2669 -1157
rect -2635 -1191 -2601 -1157
rect -2567 -1191 -2533 -1157
rect -2499 -1191 -2465 -1157
rect -2431 -1191 -2397 -1157
rect -2363 -1191 -2329 -1157
rect -2295 -1191 -2261 -1157
rect -2227 -1191 -2193 -1157
rect -2159 -1191 -2125 -1157
rect -2091 -1191 -2057 -1157
rect -2023 -1191 -1989 -1157
rect -1955 -1191 -1921 -1157
rect -1887 -1191 -1853 -1157
rect -1819 -1191 -1785 -1157
rect -1751 -1191 -1717 -1157
rect -1683 -1191 -1649 -1157
rect -1615 -1191 -1581 -1157
rect -1547 -1191 -1513 -1157
rect -1479 -1191 -1445 -1157
rect -1411 -1191 -1377 -1157
rect -1343 -1191 -1309 -1157
rect -1275 -1191 -1241 -1157
rect -1207 -1191 -1173 -1157
rect -1139 -1191 -1105 -1157
rect -1071 -1191 -1037 -1157
rect -1003 -1191 -969 -1157
rect -935 -1191 -901 -1157
rect -867 -1191 -833 -1157
rect -799 -1191 -765 -1157
rect -731 -1191 -697 -1157
rect -663 -1191 -629 -1157
rect -595 -1191 -561 -1157
rect -527 -1191 -493 -1157
rect -459 -1191 -425 -1157
rect -391 -1191 -357 -1157
rect -323 -1191 -289 -1157
rect -255 -1191 -221 -1157
rect -187 -1191 -153 -1157
rect -119 -1191 -85 -1157
rect -51 -1191 -17 -1157
rect 17 -1191 51 -1157
rect 85 -1191 119 -1157
rect 153 -1191 187 -1157
rect 221 -1191 255 -1157
rect 289 -1191 323 -1157
rect 357 -1191 391 -1157
rect 425 -1191 459 -1157
rect 493 -1191 527 -1157
rect 561 -1191 595 -1157
rect 629 -1191 663 -1157
rect 697 -1191 731 -1157
rect 765 -1191 799 -1157
rect 833 -1191 867 -1157
rect 901 -1191 935 -1157
rect 969 -1191 1003 -1157
rect 1037 -1191 1071 -1157
rect 1105 -1191 1139 -1157
rect 1173 -1191 1207 -1157
rect 1241 -1191 1275 -1157
rect 1309 -1191 1343 -1157
rect 1377 -1191 1411 -1157
rect 1445 -1191 1479 -1157
rect 1513 -1191 1547 -1157
rect 1581 -1191 1615 -1157
rect 1649 -1191 1683 -1157
rect 1717 -1191 1751 -1157
rect 1785 -1191 1819 -1157
rect 1853 -1191 1887 -1157
rect 1921 -1191 1955 -1157
rect 1989 -1191 2023 -1157
rect 2057 -1191 2091 -1157
rect 2125 -1191 2159 -1157
rect 2193 -1191 2227 -1157
rect 2261 -1191 2295 -1157
rect 2329 -1191 2363 -1157
rect 2397 -1191 2431 -1157
rect 2465 -1191 2499 -1157
rect 2533 -1191 2567 -1157
rect 2601 -1191 2635 -1157
rect 2669 -1191 2703 -1157
rect 2737 -1191 2771 -1157
rect 2805 -1191 2839 -1157
rect 2873 -1191 2907 -1157
rect 2941 -1191 2975 -1157
rect 3009 -1191 3043 -1157
rect 3077 -1191 3111 -1157
rect 3145 -1191 3179 -1157
rect 3213 -1191 3311 -1157
<< viali >>
rect -3098 1019 -3064 1053
rect -2940 1019 -2906 1053
rect -2782 1019 -2748 1053
rect -2624 1019 -2590 1053
rect -2466 1019 -2432 1053
rect -2308 1019 -2274 1053
rect -2150 1019 -2116 1053
rect -1992 1019 -1958 1053
rect -1834 1019 -1800 1053
rect -1676 1019 -1642 1053
rect -1518 1019 -1484 1053
rect -1360 1019 -1326 1053
rect -1202 1019 -1168 1053
rect -1044 1019 -1010 1053
rect -886 1019 -852 1053
rect -728 1019 -694 1053
rect -570 1019 -536 1053
rect -412 1019 -378 1053
rect -254 1019 -220 1053
rect -96 1019 -62 1053
rect 62 1019 96 1053
rect 220 1019 254 1053
rect 378 1019 412 1053
rect 536 1019 570 1053
rect 694 1019 728 1053
rect 852 1019 886 1053
rect 1010 1019 1044 1053
rect 1168 1019 1202 1053
rect 1326 1019 1360 1053
rect 1484 1019 1518 1053
rect 1642 1019 1676 1053
rect 1800 1019 1834 1053
rect 1958 1019 1992 1053
rect 2116 1019 2150 1053
rect 2274 1019 2308 1053
rect 2432 1019 2466 1053
rect 2590 1019 2624 1053
rect 2748 1019 2782 1053
rect 2906 1019 2940 1053
rect 3064 1019 3098 1053
rect -3177 923 -3143 925
rect -3177 891 -3143 923
rect -3177 821 -3143 853
rect -3177 819 -3143 821
rect -3019 923 -2985 925
rect -3019 891 -2985 923
rect -3019 821 -2985 853
rect -3019 819 -2985 821
rect -2861 923 -2827 925
rect -2861 891 -2827 923
rect -2861 821 -2827 853
rect -2861 819 -2827 821
rect -2703 923 -2669 925
rect -2703 891 -2669 923
rect -2703 821 -2669 853
rect -2703 819 -2669 821
rect -2545 923 -2511 925
rect -2545 891 -2511 923
rect -2545 821 -2511 853
rect -2545 819 -2511 821
rect -2387 923 -2353 925
rect -2387 891 -2353 923
rect -2387 821 -2353 853
rect -2387 819 -2353 821
rect -2229 923 -2195 925
rect -2229 891 -2195 923
rect -2229 821 -2195 853
rect -2229 819 -2195 821
rect -2071 923 -2037 925
rect -2071 891 -2037 923
rect -2071 821 -2037 853
rect -2071 819 -2037 821
rect -1913 923 -1879 925
rect -1913 891 -1879 923
rect -1913 821 -1879 853
rect -1913 819 -1879 821
rect -1755 923 -1721 925
rect -1755 891 -1721 923
rect -1755 821 -1721 853
rect -1755 819 -1721 821
rect -1597 923 -1563 925
rect -1597 891 -1563 923
rect -1597 821 -1563 853
rect -1597 819 -1563 821
rect -1439 923 -1405 925
rect -1439 891 -1405 923
rect -1439 821 -1405 853
rect -1439 819 -1405 821
rect -1281 923 -1247 925
rect -1281 891 -1247 923
rect -1281 821 -1247 853
rect -1281 819 -1247 821
rect -1123 923 -1089 925
rect -1123 891 -1089 923
rect -1123 821 -1089 853
rect -1123 819 -1089 821
rect -965 923 -931 925
rect -965 891 -931 923
rect -965 821 -931 853
rect -965 819 -931 821
rect -807 923 -773 925
rect -807 891 -773 923
rect -807 821 -773 853
rect -807 819 -773 821
rect -649 923 -615 925
rect -649 891 -615 923
rect -649 821 -615 853
rect -649 819 -615 821
rect -491 923 -457 925
rect -491 891 -457 923
rect -491 821 -457 853
rect -491 819 -457 821
rect -333 923 -299 925
rect -333 891 -299 923
rect -333 821 -299 853
rect -333 819 -299 821
rect -175 923 -141 925
rect -175 891 -141 923
rect -175 821 -141 853
rect -175 819 -141 821
rect -17 923 17 925
rect -17 891 17 923
rect -17 821 17 853
rect -17 819 17 821
rect 141 923 175 925
rect 141 891 175 923
rect 141 821 175 853
rect 141 819 175 821
rect 299 923 333 925
rect 299 891 333 923
rect 299 821 333 853
rect 299 819 333 821
rect 457 923 491 925
rect 457 891 491 923
rect 457 821 491 853
rect 457 819 491 821
rect 615 923 649 925
rect 615 891 649 923
rect 615 821 649 853
rect 615 819 649 821
rect 773 923 807 925
rect 773 891 807 923
rect 773 821 807 853
rect 773 819 807 821
rect 931 923 965 925
rect 931 891 965 923
rect 931 821 965 853
rect 931 819 965 821
rect 1089 923 1123 925
rect 1089 891 1123 923
rect 1089 821 1123 853
rect 1089 819 1123 821
rect 1247 923 1281 925
rect 1247 891 1281 923
rect 1247 821 1281 853
rect 1247 819 1281 821
rect 1405 923 1439 925
rect 1405 891 1439 923
rect 1405 821 1439 853
rect 1405 819 1439 821
rect 1563 923 1597 925
rect 1563 891 1597 923
rect 1563 821 1597 853
rect 1563 819 1597 821
rect 1721 923 1755 925
rect 1721 891 1755 923
rect 1721 821 1755 853
rect 1721 819 1755 821
rect 1879 923 1913 925
rect 1879 891 1913 923
rect 1879 821 1913 853
rect 1879 819 1913 821
rect 2037 923 2071 925
rect 2037 891 2071 923
rect 2037 821 2071 853
rect 2037 819 2071 821
rect 2195 923 2229 925
rect 2195 891 2229 923
rect 2195 821 2229 853
rect 2195 819 2229 821
rect 2353 923 2387 925
rect 2353 891 2387 923
rect 2353 821 2387 853
rect 2353 819 2387 821
rect 2511 923 2545 925
rect 2511 891 2545 923
rect 2511 821 2545 853
rect 2511 819 2545 821
rect 2669 923 2703 925
rect 2669 891 2703 923
rect 2669 821 2703 853
rect 2669 819 2703 821
rect 2827 923 2861 925
rect 2827 891 2861 923
rect 2827 821 2861 853
rect 2827 819 2861 821
rect 2985 923 3019 925
rect 2985 891 3019 923
rect 2985 821 3019 853
rect 2985 819 3019 821
rect 3143 923 3177 925
rect 3143 891 3177 923
rect 3143 821 3177 853
rect 3143 819 3177 821
rect -3098 691 -3064 725
rect -2940 691 -2906 725
rect -2782 691 -2748 725
rect -2624 691 -2590 725
rect -2466 691 -2432 725
rect -2308 691 -2274 725
rect -2150 691 -2116 725
rect -1992 691 -1958 725
rect -1834 691 -1800 725
rect -1676 691 -1642 725
rect -1518 691 -1484 725
rect -1360 691 -1326 725
rect -1202 691 -1168 725
rect -1044 691 -1010 725
rect -886 691 -852 725
rect -728 691 -694 725
rect -570 691 -536 725
rect -412 691 -378 725
rect -254 691 -220 725
rect -96 691 -62 725
rect 62 691 96 725
rect 220 691 254 725
rect 378 691 412 725
rect 536 691 570 725
rect 694 691 728 725
rect 852 691 886 725
rect 1010 691 1044 725
rect 1168 691 1202 725
rect 1326 691 1360 725
rect 1484 691 1518 725
rect 1642 691 1676 725
rect 1800 691 1834 725
rect 1958 691 1992 725
rect 2116 691 2150 725
rect 2274 691 2308 725
rect 2432 691 2466 725
rect 2590 691 2624 725
rect 2748 691 2782 725
rect 2906 691 2940 725
rect 3064 691 3098 725
rect -3098 583 -3064 617
rect -2940 583 -2906 617
rect -2782 583 -2748 617
rect -2624 583 -2590 617
rect -2466 583 -2432 617
rect -2308 583 -2274 617
rect -2150 583 -2116 617
rect -1992 583 -1958 617
rect -1834 583 -1800 617
rect -1676 583 -1642 617
rect -1518 583 -1484 617
rect -1360 583 -1326 617
rect -1202 583 -1168 617
rect -1044 583 -1010 617
rect -886 583 -852 617
rect -728 583 -694 617
rect -570 583 -536 617
rect -412 583 -378 617
rect -254 583 -220 617
rect -96 583 -62 617
rect 62 583 96 617
rect 220 583 254 617
rect 378 583 412 617
rect 536 583 570 617
rect 694 583 728 617
rect 852 583 886 617
rect 1010 583 1044 617
rect 1168 583 1202 617
rect 1326 583 1360 617
rect 1484 583 1518 617
rect 1642 583 1676 617
rect 1800 583 1834 617
rect 1958 583 1992 617
rect 2116 583 2150 617
rect 2274 583 2308 617
rect 2432 583 2466 617
rect 2590 583 2624 617
rect 2748 583 2782 617
rect 2906 583 2940 617
rect 3064 583 3098 617
rect -3177 487 -3143 489
rect -3177 455 -3143 487
rect -3177 385 -3143 417
rect -3177 383 -3143 385
rect -3019 487 -2985 489
rect -3019 455 -2985 487
rect -3019 385 -2985 417
rect -3019 383 -2985 385
rect -2861 487 -2827 489
rect -2861 455 -2827 487
rect -2861 385 -2827 417
rect -2861 383 -2827 385
rect -2703 487 -2669 489
rect -2703 455 -2669 487
rect -2703 385 -2669 417
rect -2703 383 -2669 385
rect -2545 487 -2511 489
rect -2545 455 -2511 487
rect -2545 385 -2511 417
rect -2545 383 -2511 385
rect -2387 487 -2353 489
rect -2387 455 -2353 487
rect -2387 385 -2353 417
rect -2387 383 -2353 385
rect -2229 487 -2195 489
rect -2229 455 -2195 487
rect -2229 385 -2195 417
rect -2229 383 -2195 385
rect -2071 487 -2037 489
rect -2071 455 -2037 487
rect -2071 385 -2037 417
rect -2071 383 -2037 385
rect -1913 487 -1879 489
rect -1913 455 -1879 487
rect -1913 385 -1879 417
rect -1913 383 -1879 385
rect -1755 487 -1721 489
rect -1755 455 -1721 487
rect -1755 385 -1721 417
rect -1755 383 -1721 385
rect -1597 487 -1563 489
rect -1597 455 -1563 487
rect -1597 385 -1563 417
rect -1597 383 -1563 385
rect -1439 487 -1405 489
rect -1439 455 -1405 487
rect -1439 385 -1405 417
rect -1439 383 -1405 385
rect -1281 487 -1247 489
rect -1281 455 -1247 487
rect -1281 385 -1247 417
rect -1281 383 -1247 385
rect -1123 487 -1089 489
rect -1123 455 -1089 487
rect -1123 385 -1089 417
rect -1123 383 -1089 385
rect -965 487 -931 489
rect -965 455 -931 487
rect -965 385 -931 417
rect -965 383 -931 385
rect -807 487 -773 489
rect -807 455 -773 487
rect -807 385 -773 417
rect -807 383 -773 385
rect -649 487 -615 489
rect -649 455 -615 487
rect -649 385 -615 417
rect -649 383 -615 385
rect -491 487 -457 489
rect -491 455 -457 487
rect -491 385 -457 417
rect -491 383 -457 385
rect -333 487 -299 489
rect -333 455 -299 487
rect -333 385 -299 417
rect -333 383 -299 385
rect -175 487 -141 489
rect -175 455 -141 487
rect -175 385 -141 417
rect -175 383 -141 385
rect -17 487 17 489
rect -17 455 17 487
rect -17 385 17 417
rect -17 383 17 385
rect 141 487 175 489
rect 141 455 175 487
rect 141 385 175 417
rect 141 383 175 385
rect 299 487 333 489
rect 299 455 333 487
rect 299 385 333 417
rect 299 383 333 385
rect 457 487 491 489
rect 457 455 491 487
rect 457 385 491 417
rect 457 383 491 385
rect 615 487 649 489
rect 615 455 649 487
rect 615 385 649 417
rect 615 383 649 385
rect 773 487 807 489
rect 773 455 807 487
rect 773 385 807 417
rect 773 383 807 385
rect 931 487 965 489
rect 931 455 965 487
rect 931 385 965 417
rect 931 383 965 385
rect 1089 487 1123 489
rect 1089 455 1123 487
rect 1089 385 1123 417
rect 1089 383 1123 385
rect 1247 487 1281 489
rect 1247 455 1281 487
rect 1247 385 1281 417
rect 1247 383 1281 385
rect 1405 487 1439 489
rect 1405 455 1439 487
rect 1405 385 1439 417
rect 1405 383 1439 385
rect 1563 487 1597 489
rect 1563 455 1597 487
rect 1563 385 1597 417
rect 1563 383 1597 385
rect 1721 487 1755 489
rect 1721 455 1755 487
rect 1721 385 1755 417
rect 1721 383 1755 385
rect 1879 487 1913 489
rect 1879 455 1913 487
rect 1879 385 1913 417
rect 1879 383 1913 385
rect 2037 487 2071 489
rect 2037 455 2071 487
rect 2037 385 2071 417
rect 2037 383 2071 385
rect 2195 487 2229 489
rect 2195 455 2229 487
rect 2195 385 2229 417
rect 2195 383 2229 385
rect 2353 487 2387 489
rect 2353 455 2387 487
rect 2353 385 2387 417
rect 2353 383 2387 385
rect 2511 487 2545 489
rect 2511 455 2545 487
rect 2511 385 2545 417
rect 2511 383 2545 385
rect 2669 487 2703 489
rect 2669 455 2703 487
rect 2669 385 2703 417
rect 2669 383 2703 385
rect 2827 487 2861 489
rect 2827 455 2861 487
rect 2827 385 2861 417
rect 2827 383 2861 385
rect 2985 487 3019 489
rect 2985 455 3019 487
rect 2985 385 3019 417
rect 2985 383 3019 385
rect 3143 487 3177 489
rect 3143 455 3177 487
rect 3143 385 3177 417
rect 3143 383 3177 385
rect -3098 255 -3064 289
rect -2940 255 -2906 289
rect -2782 255 -2748 289
rect -2624 255 -2590 289
rect -2466 255 -2432 289
rect -2308 255 -2274 289
rect -2150 255 -2116 289
rect -1992 255 -1958 289
rect -1834 255 -1800 289
rect -1676 255 -1642 289
rect -1518 255 -1484 289
rect -1360 255 -1326 289
rect -1202 255 -1168 289
rect -1044 255 -1010 289
rect -886 255 -852 289
rect -728 255 -694 289
rect -570 255 -536 289
rect -412 255 -378 289
rect -254 255 -220 289
rect -96 255 -62 289
rect 62 255 96 289
rect 220 255 254 289
rect 378 255 412 289
rect 536 255 570 289
rect 694 255 728 289
rect 852 255 886 289
rect 1010 255 1044 289
rect 1168 255 1202 289
rect 1326 255 1360 289
rect 1484 255 1518 289
rect 1642 255 1676 289
rect 1800 255 1834 289
rect 1958 255 1992 289
rect 2116 255 2150 289
rect 2274 255 2308 289
rect 2432 255 2466 289
rect 2590 255 2624 289
rect 2748 255 2782 289
rect 2906 255 2940 289
rect 3064 255 3098 289
rect -3098 147 -3064 181
rect -2940 147 -2906 181
rect -2782 147 -2748 181
rect -2624 147 -2590 181
rect -2466 147 -2432 181
rect -2308 147 -2274 181
rect -2150 147 -2116 181
rect -1992 147 -1958 181
rect -1834 147 -1800 181
rect -1676 147 -1642 181
rect -1518 147 -1484 181
rect -1360 147 -1326 181
rect -1202 147 -1168 181
rect -1044 147 -1010 181
rect -886 147 -852 181
rect -728 147 -694 181
rect -570 147 -536 181
rect -412 147 -378 181
rect -254 147 -220 181
rect -96 147 -62 181
rect 62 147 96 181
rect 220 147 254 181
rect 378 147 412 181
rect 536 147 570 181
rect 694 147 728 181
rect 852 147 886 181
rect 1010 147 1044 181
rect 1168 147 1202 181
rect 1326 147 1360 181
rect 1484 147 1518 181
rect 1642 147 1676 181
rect 1800 147 1834 181
rect 1958 147 1992 181
rect 2116 147 2150 181
rect 2274 147 2308 181
rect 2432 147 2466 181
rect 2590 147 2624 181
rect 2748 147 2782 181
rect 2906 147 2940 181
rect 3064 147 3098 181
rect -3177 51 -3143 53
rect -3177 19 -3143 51
rect -3177 -51 -3143 -19
rect -3177 -53 -3143 -51
rect -3019 51 -2985 53
rect -3019 19 -2985 51
rect -3019 -51 -2985 -19
rect -3019 -53 -2985 -51
rect -2861 51 -2827 53
rect -2861 19 -2827 51
rect -2861 -51 -2827 -19
rect -2861 -53 -2827 -51
rect -2703 51 -2669 53
rect -2703 19 -2669 51
rect -2703 -51 -2669 -19
rect -2703 -53 -2669 -51
rect -2545 51 -2511 53
rect -2545 19 -2511 51
rect -2545 -51 -2511 -19
rect -2545 -53 -2511 -51
rect -2387 51 -2353 53
rect -2387 19 -2353 51
rect -2387 -51 -2353 -19
rect -2387 -53 -2353 -51
rect -2229 51 -2195 53
rect -2229 19 -2195 51
rect -2229 -51 -2195 -19
rect -2229 -53 -2195 -51
rect -2071 51 -2037 53
rect -2071 19 -2037 51
rect -2071 -51 -2037 -19
rect -2071 -53 -2037 -51
rect -1913 51 -1879 53
rect -1913 19 -1879 51
rect -1913 -51 -1879 -19
rect -1913 -53 -1879 -51
rect -1755 51 -1721 53
rect -1755 19 -1721 51
rect -1755 -51 -1721 -19
rect -1755 -53 -1721 -51
rect -1597 51 -1563 53
rect -1597 19 -1563 51
rect -1597 -51 -1563 -19
rect -1597 -53 -1563 -51
rect -1439 51 -1405 53
rect -1439 19 -1405 51
rect -1439 -51 -1405 -19
rect -1439 -53 -1405 -51
rect -1281 51 -1247 53
rect -1281 19 -1247 51
rect -1281 -51 -1247 -19
rect -1281 -53 -1247 -51
rect -1123 51 -1089 53
rect -1123 19 -1089 51
rect -1123 -51 -1089 -19
rect -1123 -53 -1089 -51
rect -965 51 -931 53
rect -965 19 -931 51
rect -965 -51 -931 -19
rect -965 -53 -931 -51
rect -807 51 -773 53
rect -807 19 -773 51
rect -807 -51 -773 -19
rect -807 -53 -773 -51
rect -649 51 -615 53
rect -649 19 -615 51
rect -649 -51 -615 -19
rect -649 -53 -615 -51
rect -491 51 -457 53
rect -491 19 -457 51
rect -491 -51 -457 -19
rect -491 -53 -457 -51
rect -333 51 -299 53
rect -333 19 -299 51
rect -333 -51 -299 -19
rect -333 -53 -299 -51
rect -175 51 -141 53
rect -175 19 -141 51
rect -175 -51 -141 -19
rect -175 -53 -141 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 141 51 175 53
rect 141 19 175 51
rect 141 -51 175 -19
rect 141 -53 175 -51
rect 299 51 333 53
rect 299 19 333 51
rect 299 -51 333 -19
rect 299 -53 333 -51
rect 457 51 491 53
rect 457 19 491 51
rect 457 -51 491 -19
rect 457 -53 491 -51
rect 615 51 649 53
rect 615 19 649 51
rect 615 -51 649 -19
rect 615 -53 649 -51
rect 773 51 807 53
rect 773 19 807 51
rect 773 -51 807 -19
rect 773 -53 807 -51
rect 931 51 965 53
rect 931 19 965 51
rect 931 -51 965 -19
rect 931 -53 965 -51
rect 1089 51 1123 53
rect 1089 19 1123 51
rect 1089 -51 1123 -19
rect 1089 -53 1123 -51
rect 1247 51 1281 53
rect 1247 19 1281 51
rect 1247 -51 1281 -19
rect 1247 -53 1281 -51
rect 1405 51 1439 53
rect 1405 19 1439 51
rect 1405 -51 1439 -19
rect 1405 -53 1439 -51
rect 1563 51 1597 53
rect 1563 19 1597 51
rect 1563 -51 1597 -19
rect 1563 -53 1597 -51
rect 1721 51 1755 53
rect 1721 19 1755 51
rect 1721 -51 1755 -19
rect 1721 -53 1755 -51
rect 1879 51 1913 53
rect 1879 19 1913 51
rect 1879 -51 1913 -19
rect 1879 -53 1913 -51
rect 2037 51 2071 53
rect 2037 19 2071 51
rect 2037 -51 2071 -19
rect 2037 -53 2071 -51
rect 2195 51 2229 53
rect 2195 19 2229 51
rect 2195 -51 2229 -19
rect 2195 -53 2229 -51
rect 2353 51 2387 53
rect 2353 19 2387 51
rect 2353 -51 2387 -19
rect 2353 -53 2387 -51
rect 2511 51 2545 53
rect 2511 19 2545 51
rect 2511 -51 2545 -19
rect 2511 -53 2545 -51
rect 2669 51 2703 53
rect 2669 19 2703 51
rect 2669 -51 2703 -19
rect 2669 -53 2703 -51
rect 2827 51 2861 53
rect 2827 19 2861 51
rect 2827 -51 2861 -19
rect 2827 -53 2861 -51
rect 2985 51 3019 53
rect 2985 19 3019 51
rect 2985 -51 3019 -19
rect 2985 -53 3019 -51
rect 3143 51 3177 53
rect 3143 19 3177 51
rect 3143 -51 3177 -19
rect 3143 -53 3177 -51
rect -3098 -181 -3064 -147
rect -2940 -181 -2906 -147
rect -2782 -181 -2748 -147
rect -2624 -181 -2590 -147
rect -2466 -181 -2432 -147
rect -2308 -181 -2274 -147
rect -2150 -181 -2116 -147
rect -1992 -181 -1958 -147
rect -1834 -181 -1800 -147
rect -1676 -181 -1642 -147
rect -1518 -181 -1484 -147
rect -1360 -181 -1326 -147
rect -1202 -181 -1168 -147
rect -1044 -181 -1010 -147
rect -886 -181 -852 -147
rect -728 -181 -694 -147
rect -570 -181 -536 -147
rect -412 -181 -378 -147
rect -254 -181 -220 -147
rect -96 -181 -62 -147
rect 62 -181 96 -147
rect 220 -181 254 -147
rect 378 -181 412 -147
rect 536 -181 570 -147
rect 694 -181 728 -147
rect 852 -181 886 -147
rect 1010 -181 1044 -147
rect 1168 -181 1202 -147
rect 1326 -181 1360 -147
rect 1484 -181 1518 -147
rect 1642 -181 1676 -147
rect 1800 -181 1834 -147
rect 1958 -181 1992 -147
rect 2116 -181 2150 -147
rect 2274 -181 2308 -147
rect 2432 -181 2466 -147
rect 2590 -181 2624 -147
rect 2748 -181 2782 -147
rect 2906 -181 2940 -147
rect 3064 -181 3098 -147
rect -3098 -289 -3064 -255
rect -2940 -289 -2906 -255
rect -2782 -289 -2748 -255
rect -2624 -289 -2590 -255
rect -2466 -289 -2432 -255
rect -2308 -289 -2274 -255
rect -2150 -289 -2116 -255
rect -1992 -289 -1958 -255
rect -1834 -289 -1800 -255
rect -1676 -289 -1642 -255
rect -1518 -289 -1484 -255
rect -1360 -289 -1326 -255
rect -1202 -289 -1168 -255
rect -1044 -289 -1010 -255
rect -886 -289 -852 -255
rect -728 -289 -694 -255
rect -570 -289 -536 -255
rect -412 -289 -378 -255
rect -254 -289 -220 -255
rect -96 -289 -62 -255
rect 62 -289 96 -255
rect 220 -289 254 -255
rect 378 -289 412 -255
rect 536 -289 570 -255
rect 694 -289 728 -255
rect 852 -289 886 -255
rect 1010 -289 1044 -255
rect 1168 -289 1202 -255
rect 1326 -289 1360 -255
rect 1484 -289 1518 -255
rect 1642 -289 1676 -255
rect 1800 -289 1834 -255
rect 1958 -289 1992 -255
rect 2116 -289 2150 -255
rect 2274 -289 2308 -255
rect 2432 -289 2466 -255
rect 2590 -289 2624 -255
rect 2748 -289 2782 -255
rect 2906 -289 2940 -255
rect 3064 -289 3098 -255
rect -3177 -385 -3143 -383
rect -3177 -417 -3143 -385
rect -3177 -487 -3143 -455
rect -3177 -489 -3143 -487
rect -3019 -385 -2985 -383
rect -3019 -417 -2985 -385
rect -3019 -487 -2985 -455
rect -3019 -489 -2985 -487
rect -2861 -385 -2827 -383
rect -2861 -417 -2827 -385
rect -2861 -487 -2827 -455
rect -2861 -489 -2827 -487
rect -2703 -385 -2669 -383
rect -2703 -417 -2669 -385
rect -2703 -487 -2669 -455
rect -2703 -489 -2669 -487
rect -2545 -385 -2511 -383
rect -2545 -417 -2511 -385
rect -2545 -487 -2511 -455
rect -2545 -489 -2511 -487
rect -2387 -385 -2353 -383
rect -2387 -417 -2353 -385
rect -2387 -487 -2353 -455
rect -2387 -489 -2353 -487
rect -2229 -385 -2195 -383
rect -2229 -417 -2195 -385
rect -2229 -487 -2195 -455
rect -2229 -489 -2195 -487
rect -2071 -385 -2037 -383
rect -2071 -417 -2037 -385
rect -2071 -487 -2037 -455
rect -2071 -489 -2037 -487
rect -1913 -385 -1879 -383
rect -1913 -417 -1879 -385
rect -1913 -487 -1879 -455
rect -1913 -489 -1879 -487
rect -1755 -385 -1721 -383
rect -1755 -417 -1721 -385
rect -1755 -487 -1721 -455
rect -1755 -489 -1721 -487
rect -1597 -385 -1563 -383
rect -1597 -417 -1563 -385
rect -1597 -487 -1563 -455
rect -1597 -489 -1563 -487
rect -1439 -385 -1405 -383
rect -1439 -417 -1405 -385
rect -1439 -487 -1405 -455
rect -1439 -489 -1405 -487
rect -1281 -385 -1247 -383
rect -1281 -417 -1247 -385
rect -1281 -487 -1247 -455
rect -1281 -489 -1247 -487
rect -1123 -385 -1089 -383
rect -1123 -417 -1089 -385
rect -1123 -487 -1089 -455
rect -1123 -489 -1089 -487
rect -965 -385 -931 -383
rect -965 -417 -931 -385
rect -965 -487 -931 -455
rect -965 -489 -931 -487
rect -807 -385 -773 -383
rect -807 -417 -773 -385
rect -807 -487 -773 -455
rect -807 -489 -773 -487
rect -649 -385 -615 -383
rect -649 -417 -615 -385
rect -649 -487 -615 -455
rect -649 -489 -615 -487
rect -491 -385 -457 -383
rect -491 -417 -457 -385
rect -491 -487 -457 -455
rect -491 -489 -457 -487
rect -333 -385 -299 -383
rect -333 -417 -299 -385
rect -333 -487 -299 -455
rect -333 -489 -299 -487
rect -175 -385 -141 -383
rect -175 -417 -141 -385
rect -175 -487 -141 -455
rect -175 -489 -141 -487
rect -17 -385 17 -383
rect -17 -417 17 -385
rect -17 -487 17 -455
rect -17 -489 17 -487
rect 141 -385 175 -383
rect 141 -417 175 -385
rect 141 -487 175 -455
rect 141 -489 175 -487
rect 299 -385 333 -383
rect 299 -417 333 -385
rect 299 -487 333 -455
rect 299 -489 333 -487
rect 457 -385 491 -383
rect 457 -417 491 -385
rect 457 -487 491 -455
rect 457 -489 491 -487
rect 615 -385 649 -383
rect 615 -417 649 -385
rect 615 -487 649 -455
rect 615 -489 649 -487
rect 773 -385 807 -383
rect 773 -417 807 -385
rect 773 -487 807 -455
rect 773 -489 807 -487
rect 931 -385 965 -383
rect 931 -417 965 -385
rect 931 -487 965 -455
rect 931 -489 965 -487
rect 1089 -385 1123 -383
rect 1089 -417 1123 -385
rect 1089 -487 1123 -455
rect 1089 -489 1123 -487
rect 1247 -385 1281 -383
rect 1247 -417 1281 -385
rect 1247 -487 1281 -455
rect 1247 -489 1281 -487
rect 1405 -385 1439 -383
rect 1405 -417 1439 -385
rect 1405 -487 1439 -455
rect 1405 -489 1439 -487
rect 1563 -385 1597 -383
rect 1563 -417 1597 -385
rect 1563 -487 1597 -455
rect 1563 -489 1597 -487
rect 1721 -385 1755 -383
rect 1721 -417 1755 -385
rect 1721 -487 1755 -455
rect 1721 -489 1755 -487
rect 1879 -385 1913 -383
rect 1879 -417 1913 -385
rect 1879 -487 1913 -455
rect 1879 -489 1913 -487
rect 2037 -385 2071 -383
rect 2037 -417 2071 -385
rect 2037 -487 2071 -455
rect 2037 -489 2071 -487
rect 2195 -385 2229 -383
rect 2195 -417 2229 -385
rect 2195 -487 2229 -455
rect 2195 -489 2229 -487
rect 2353 -385 2387 -383
rect 2353 -417 2387 -385
rect 2353 -487 2387 -455
rect 2353 -489 2387 -487
rect 2511 -385 2545 -383
rect 2511 -417 2545 -385
rect 2511 -487 2545 -455
rect 2511 -489 2545 -487
rect 2669 -385 2703 -383
rect 2669 -417 2703 -385
rect 2669 -487 2703 -455
rect 2669 -489 2703 -487
rect 2827 -385 2861 -383
rect 2827 -417 2861 -385
rect 2827 -487 2861 -455
rect 2827 -489 2861 -487
rect 2985 -385 3019 -383
rect 2985 -417 3019 -385
rect 2985 -487 3019 -455
rect 2985 -489 3019 -487
rect 3143 -385 3177 -383
rect 3143 -417 3177 -385
rect 3143 -487 3177 -455
rect 3143 -489 3177 -487
rect -3098 -617 -3064 -583
rect -2940 -617 -2906 -583
rect -2782 -617 -2748 -583
rect -2624 -617 -2590 -583
rect -2466 -617 -2432 -583
rect -2308 -617 -2274 -583
rect -2150 -617 -2116 -583
rect -1992 -617 -1958 -583
rect -1834 -617 -1800 -583
rect -1676 -617 -1642 -583
rect -1518 -617 -1484 -583
rect -1360 -617 -1326 -583
rect -1202 -617 -1168 -583
rect -1044 -617 -1010 -583
rect -886 -617 -852 -583
rect -728 -617 -694 -583
rect -570 -617 -536 -583
rect -412 -617 -378 -583
rect -254 -617 -220 -583
rect -96 -617 -62 -583
rect 62 -617 96 -583
rect 220 -617 254 -583
rect 378 -617 412 -583
rect 536 -617 570 -583
rect 694 -617 728 -583
rect 852 -617 886 -583
rect 1010 -617 1044 -583
rect 1168 -617 1202 -583
rect 1326 -617 1360 -583
rect 1484 -617 1518 -583
rect 1642 -617 1676 -583
rect 1800 -617 1834 -583
rect 1958 -617 1992 -583
rect 2116 -617 2150 -583
rect 2274 -617 2308 -583
rect 2432 -617 2466 -583
rect 2590 -617 2624 -583
rect 2748 -617 2782 -583
rect 2906 -617 2940 -583
rect 3064 -617 3098 -583
rect -3098 -725 -3064 -691
rect -2940 -725 -2906 -691
rect -2782 -725 -2748 -691
rect -2624 -725 -2590 -691
rect -2466 -725 -2432 -691
rect -2308 -725 -2274 -691
rect -2150 -725 -2116 -691
rect -1992 -725 -1958 -691
rect -1834 -725 -1800 -691
rect -1676 -725 -1642 -691
rect -1518 -725 -1484 -691
rect -1360 -725 -1326 -691
rect -1202 -725 -1168 -691
rect -1044 -725 -1010 -691
rect -886 -725 -852 -691
rect -728 -725 -694 -691
rect -570 -725 -536 -691
rect -412 -725 -378 -691
rect -254 -725 -220 -691
rect -96 -725 -62 -691
rect 62 -725 96 -691
rect 220 -725 254 -691
rect 378 -725 412 -691
rect 536 -725 570 -691
rect 694 -725 728 -691
rect 852 -725 886 -691
rect 1010 -725 1044 -691
rect 1168 -725 1202 -691
rect 1326 -725 1360 -691
rect 1484 -725 1518 -691
rect 1642 -725 1676 -691
rect 1800 -725 1834 -691
rect 1958 -725 1992 -691
rect 2116 -725 2150 -691
rect 2274 -725 2308 -691
rect 2432 -725 2466 -691
rect 2590 -725 2624 -691
rect 2748 -725 2782 -691
rect 2906 -725 2940 -691
rect 3064 -725 3098 -691
rect -3177 -821 -3143 -819
rect -3177 -853 -3143 -821
rect -3177 -923 -3143 -891
rect -3177 -925 -3143 -923
rect -3019 -821 -2985 -819
rect -3019 -853 -2985 -821
rect -3019 -923 -2985 -891
rect -3019 -925 -2985 -923
rect -2861 -821 -2827 -819
rect -2861 -853 -2827 -821
rect -2861 -923 -2827 -891
rect -2861 -925 -2827 -923
rect -2703 -821 -2669 -819
rect -2703 -853 -2669 -821
rect -2703 -923 -2669 -891
rect -2703 -925 -2669 -923
rect -2545 -821 -2511 -819
rect -2545 -853 -2511 -821
rect -2545 -923 -2511 -891
rect -2545 -925 -2511 -923
rect -2387 -821 -2353 -819
rect -2387 -853 -2353 -821
rect -2387 -923 -2353 -891
rect -2387 -925 -2353 -923
rect -2229 -821 -2195 -819
rect -2229 -853 -2195 -821
rect -2229 -923 -2195 -891
rect -2229 -925 -2195 -923
rect -2071 -821 -2037 -819
rect -2071 -853 -2037 -821
rect -2071 -923 -2037 -891
rect -2071 -925 -2037 -923
rect -1913 -821 -1879 -819
rect -1913 -853 -1879 -821
rect -1913 -923 -1879 -891
rect -1913 -925 -1879 -923
rect -1755 -821 -1721 -819
rect -1755 -853 -1721 -821
rect -1755 -923 -1721 -891
rect -1755 -925 -1721 -923
rect -1597 -821 -1563 -819
rect -1597 -853 -1563 -821
rect -1597 -923 -1563 -891
rect -1597 -925 -1563 -923
rect -1439 -821 -1405 -819
rect -1439 -853 -1405 -821
rect -1439 -923 -1405 -891
rect -1439 -925 -1405 -923
rect -1281 -821 -1247 -819
rect -1281 -853 -1247 -821
rect -1281 -923 -1247 -891
rect -1281 -925 -1247 -923
rect -1123 -821 -1089 -819
rect -1123 -853 -1089 -821
rect -1123 -923 -1089 -891
rect -1123 -925 -1089 -923
rect -965 -821 -931 -819
rect -965 -853 -931 -821
rect -965 -923 -931 -891
rect -965 -925 -931 -923
rect -807 -821 -773 -819
rect -807 -853 -773 -821
rect -807 -923 -773 -891
rect -807 -925 -773 -923
rect -649 -821 -615 -819
rect -649 -853 -615 -821
rect -649 -923 -615 -891
rect -649 -925 -615 -923
rect -491 -821 -457 -819
rect -491 -853 -457 -821
rect -491 -923 -457 -891
rect -491 -925 -457 -923
rect -333 -821 -299 -819
rect -333 -853 -299 -821
rect -333 -923 -299 -891
rect -333 -925 -299 -923
rect -175 -821 -141 -819
rect -175 -853 -141 -821
rect -175 -923 -141 -891
rect -175 -925 -141 -923
rect -17 -821 17 -819
rect -17 -853 17 -821
rect -17 -923 17 -891
rect -17 -925 17 -923
rect 141 -821 175 -819
rect 141 -853 175 -821
rect 141 -923 175 -891
rect 141 -925 175 -923
rect 299 -821 333 -819
rect 299 -853 333 -821
rect 299 -923 333 -891
rect 299 -925 333 -923
rect 457 -821 491 -819
rect 457 -853 491 -821
rect 457 -923 491 -891
rect 457 -925 491 -923
rect 615 -821 649 -819
rect 615 -853 649 -821
rect 615 -923 649 -891
rect 615 -925 649 -923
rect 773 -821 807 -819
rect 773 -853 807 -821
rect 773 -923 807 -891
rect 773 -925 807 -923
rect 931 -821 965 -819
rect 931 -853 965 -821
rect 931 -923 965 -891
rect 931 -925 965 -923
rect 1089 -821 1123 -819
rect 1089 -853 1123 -821
rect 1089 -923 1123 -891
rect 1089 -925 1123 -923
rect 1247 -821 1281 -819
rect 1247 -853 1281 -821
rect 1247 -923 1281 -891
rect 1247 -925 1281 -923
rect 1405 -821 1439 -819
rect 1405 -853 1439 -821
rect 1405 -923 1439 -891
rect 1405 -925 1439 -923
rect 1563 -821 1597 -819
rect 1563 -853 1597 -821
rect 1563 -923 1597 -891
rect 1563 -925 1597 -923
rect 1721 -821 1755 -819
rect 1721 -853 1755 -821
rect 1721 -923 1755 -891
rect 1721 -925 1755 -923
rect 1879 -821 1913 -819
rect 1879 -853 1913 -821
rect 1879 -923 1913 -891
rect 1879 -925 1913 -923
rect 2037 -821 2071 -819
rect 2037 -853 2071 -821
rect 2037 -923 2071 -891
rect 2037 -925 2071 -923
rect 2195 -821 2229 -819
rect 2195 -853 2229 -821
rect 2195 -923 2229 -891
rect 2195 -925 2229 -923
rect 2353 -821 2387 -819
rect 2353 -853 2387 -821
rect 2353 -923 2387 -891
rect 2353 -925 2387 -923
rect 2511 -821 2545 -819
rect 2511 -853 2545 -821
rect 2511 -923 2545 -891
rect 2511 -925 2545 -923
rect 2669 -821 2703 -819
rect 2669 -853 2703 -821
rect 2669 -923 2703 -891
rect 2669 -925 2703 -923
rect 2827 -821 2861 -819
rect 2827 -853 2861 -821
rect 2827 -923 2861 -891
rect 2827 -925 2861 -923
rect 2985 -821 3019 -819
rect 2985 -853 3019 -821
rect 2985 -923 3019 -891
rect 2985 -925 3019 -923
rect 3143 -821 3177 -819
rect 3143 -853 3177 -821
rect 3143 -923 3177 -891
rect 3143 -925 3177 -923
rect -3098 -1053 -3064 -1019
rect -2940 -1053 -2906 -1019
rect -2782 -1053 -2748 -1019
rect -2624 -1053 -2590 -1019
rect -2466 -1053 -2432 -1019
rect -2308 -1053 -2274 -1019
rect -2150 -1053 -2116 -1019
rect -1992 -1053 -1958 -1019
rect -1834 -1053 -1800 -1019
rect -1676 -1053 -1642 -1019
rect -1518 -1053 -1484 -1019
rect -1360 -1053 -1326 -1019
rect -1202 -1053 -1168 -1019
rect -1044 -1053 -1010 -1019
rect -886 -1053 -852 -1019
rect -728 -1053 -694 -1019
rect -570 -1053 -536 -1019
rect -412 -1053 -378 -1019
rect -254 -1053 -220 -1019
rect -96 -1053 -62 -1019
rect 62 -1053 96 -1019
rect 220 -1053 254 -1019
rect 378 -1053 412 -1019
rect 536 -1053 570 -1019
rect 694 -1053 728 -1019
rect 852 -1053 886 -1019
rect 1010 -1053 1044 -1019
rect 1168 -1053 1202 -1019
rect 1326 -1053 1360 -1019
rect 1484 -1053 1518 -1019
rect 1642 -1053 1676 -1019
rect 1800 -1053 1834 -1019
rect 1958 -1053 1992 -1019
rect 2116 -1053 2150 -1019
rect 2274 -1053 2308 -1019
rect 2432 -1053 2466 -1019
rect 2590 -1053 2624 -1019
rect 2748 -1053 2782 -1019
rect 2906 -1053 2940 -1019
rect 3064 -1053 3098 -1019
<< metal1 >>
rect -3127 1053 -3035 1059
rect -3127 1019 -3098 1053
rect -3064 1019 -3035 1053
rect -3127 1013 -3035 1019
rect -2969 1053 -2877 1059
rect -2969 1019 -2940 1053
rect -2906 1019 -2877 1053
rect -2969 1013 -2877 1019
rect -2811 1053 -2719 1059
rect -2811 1019 -2782 1053
rect -2748 1019 -2719 1053
rect -2811 1013 -2719 1019
rect -2653 1053 -2561 1059
rect -2653 1019 -2624 1053
rect -2590 1019 -2561 1053
rect -2653 1013 -2561 1019
rect -2495 1053 -2403 1059
rect -2495 1019 -2466 1053
rect -2432 1019 -2403 1053
rect -2495 1013 -2403 1019
rect -2337 1053 -2245 1059
rect -2337 1019 -2308 1053
rect -2274 1019 -2245 1053
rect -2337 1013 -2245 1019
rect -2179 1053 -2087 1059
rect -2179 1019 -2150 1053
rect -2116 1019 -2087 1053
rect -2179 1013 -2087 1019
rect -2021 1053 -1929 1059
rect -2021 1019 -1992 1053
rect -1958 1019 -1929 1053
rect -2021 1013 -1929 1019
rect -1863 1053 -1771 1059
rect -1863 1019 -1834 1053
rect -1800 1019 -1771 1053
rect -1863 1013 -1771 1019
rect -1705 1053 -1613 1059
rect -1705 1019 -1676 1053
rect -1642 1019 -1613 1053
rect -1705 1013 -1613 1019
rect -1547 1053 -1455 1059
rect -1547 1019 -1518 1053
rect -1484 1019 -1455 1053
rect -1547 1013 -1455 1019
rect -1389 1053 -1297 1059
rect -1389 1019 -1360 1053
rect -1326 1019 -1297 1053
rect -1389 1013 -1297 1019
rect -1231 1053 -1139 1059
rect -1231 1019 -1202 1053
rect -1168 1019 -1139 1053
rect -1231 1013 -1139 1019
rect -1073 1053 -981 1059
rect -1073 1019 -1044 1053
rect -1010 1019 -981 1053
rect -1073 1013 -981 1019
rect -915 1053 -823 1059
rect -915 1019 -886 1053
rect -852 1019 -823 1053
rect -915 1013 -823 1019
rect -757 1053 -665 1059
rect -757 1019 -728 1053
rect -694 1019 -665 1053
rect -757 1013 -665 1019
rect -599 1053 -507 1059
rect -599 1019 -570 1053
rect -536 1019 -507 1053
rect -599 1013 -507 1019
rect -441 1053 -349 1059
rect -441 1019 -412 1053
rect -378 1019 -349 1053
rect -441 1013 -349 1019
rect -283 1053 -191 1059
rect -283 1019 -254 1053
rect -220 1019 -191 1053
rect -283 1013 -191 1019
rect -125 1053 -33 1059
rect -125 1019 -96 1053
rect -62 1019 -33 1053
rect -125 1013 -33 1019
rect 33 1053 125 1059
rect 33 1019 62 1053
rect 96 1019 125 1053
rect 33 1013 125 1019
rect 191 1053 283 1059
rect 191 1019 220 1053
rect 254 1019 283 1053
rect 191 1013 283 1019
rect 349 1053 441 1059
rect 349 1019 378 1053
rect 412 1019 441 1053
rect 349 1013 441 1019
rect 507 1053 599 1059
rect 507 1019 536 1053
rect 570 1019 599 1053
rect 507 1013 599 1019
rect 665 1053 757 1059
rect 665 1019 694 1053
rect 728 1019 757 1053
rect 665 1013 757 1019
rect 823 1053 915 1059
rect 823 1019 852 1053
rect 886 1019 915 1053
rect 823 1013 915 1019
rect 981 1053 1073 1059
rect 981 1019 1010 1053
rect 1044 1019 1073 1053
rect 981 1013 1073 1019
rect 1139 1053 1231 1059
rect 1139 1019 1168 1053
rect 1202 1019 1231 1053
rect 1139 1013 1231 1019
rect 1297 1053 1389 1059
rect 1297 1019 1326 1053
rect 1360 1019 1389 1053
rect 1297 1013 1389 1019
rect 1455 1053 1547 1059
rect 1455 1019 1484 1053
rect 1518 1019 1547 1053
rect 1455 1013 1547 1019
rect 1613 1053 1705 1059
rect 1613 1019 1642 1053
rect 1676 1019 1705 1053
rect 1613 1013 1705 1019
rect 1771 1053 1863 1059
rect 1771 1019 1800 1053
rect 1834 1019 1863 1053
rect 1771 1013 1863 1019
rect 1929 1053 2021 1059
rect 1929 1019 1958 1053
rect 1992 1019 2021 1053
rect 1929 1013 2021 1019
rect 2087 1053 2179 1059
rect 2087 1019 2116 1053
rect 2150 1019 2179 1053
rect 2087 1013 2179 1019
rect 2245 1053 2337 1059
rect 2245 1019 2274 1053
rect 2308 1019 2337 1053
rect 2245 1013 2337 1019
rect 2403 1053 2495 1059
rect 2403 1019 2432 1053
rect 2466 1019 2495 1053
rect 2403 1013 2495 1019
rect 2561 1053 2653 1059
rect 2561 1019 2590 1053
rect 2624 1019 2653 1053
rect 2561 1013 2653 1019
rect 2719 1053 2811 1059
rect 2719 1019 2748 1053
rect 2782 1019 2811 1053
rect 2719 1013 2811 1019
rect 2877 1053 2969 1059
rect 2877 1019 2906 1053
rect 2940 1019 2969 1053
rect 2877 1013 2969 1019
rect 3035 1053 3127 1059
rect 3035 1019 3064 1053
rect 3098 1019 3127 1053
rect 3035 1013 3127 1019
rect -3183 925 -3137 972
rect -3183 891 -3177 925
rect -3143 891 -3137 925
rect -3183 853 -3137 891
rect -3183 819 -3177 853
rect -3143 819 -3137 853
rect -3183 772 -3137 819
rect -3025 925 -2979 972
rect -3025 891 -3019 925
rect -2985 891 -2979 925
rect -3025 853 -2979 891
rect -3025 819 -3019 853
rect -2985 819 -2979 853
rect -3025 772 -2979 819
rect -2867 925 -2821 972
rect -2867 891 -2861 925
rect -2827 891 -2821 925
rect -2867 853 -2821 891
rect -2867 819 -2861 853
rect -2827 819 -2821 853
rect -2867 772 -2821 819
rect -2709 925 -2663 972
rect -2709 891 -2703 925
rect -2669 891 -2663 925
rect -2709 853 -2663 891
rect -2709 819 -2703 853
rect -2669 819 -2663 853
rect -2709 772 -2663 819
rect -2551 925 -2505 972
rect -2551 891 -2545 925
rect -2511 891 -2505 925
rect -2551 853 -2505 891
rect -2551 819 -2545 853
rect -2511 819 -2505 853
rect -2551 772 -2505 819
rect -2393 925 -2347 972
rect -2393 891 -2387 925
rect -2353 891 -2347 925
rect -2393 853 -2347 891
rect -2393 819 -2387 853
rect -2353 819 -2347 853
rect -2393 772 -2347 819
rect -2235 925 -2189 972
rect -2235 891 -2229 925
rect -2195 891 -2189 925
rect -2235 853 -2189 891
rect -2235 819 -2229 853
rect -2195 819 -2189 853
rect -2235 772 -2189 819
rect -2077 925 -2031 972
rect -2077 891 -2071 925
rect -2037 891 -2031 925
rect -2077 853 -2031 891
rect -2077 819 -2071 853
rect -2037 819 -2031 853
rect -2077 772 -2031 819
rect -1919 925 -1873 972
rect -1919 891 -1913 925
rect -1879 891 -1873 925
rect -1919 853 -1873 891
rect -1919 819 -1913 853
rect -1879 819 -1873 853
rect -1919 772 -1873 819
rect -1761 925 -1715 972
rect -1761 891 -1755 925
rect -1721 891 -1715 925
rect -1761 853 -1715 891
rect -1761 819 -1755 853
rect -1721 819 -1715 853
rect -1761 772 -1715 819
rect -1603 925 -1557 972
rect -1603 891 -1597 925
rect -1563 891 -1557 925
rect -1603 853 -1557 891
rect -1603 819 -1597 853
rect -1563 819 -1557 853
rect -1603 772 -1557 819
rect -1445 925 -1399 972
rect -1445 891 -1439 925
rect -1405 891 -1399 925
rect -1445 853 -1399 891
rect -1445 819 -1439 853
rect -1405 819 -1399 853
rect -1445 772 -1399 819
rect -1287 925 -1241 972
rect -1287 891 -1281 925
rect -1247 891 -1241 925
rect -1287 853 -1241 891
rect -1287 819 -1281 853
rect -1247 819 -1241 853
rect -1287 772 -1241 819
rect -1129 925 -1083 972
rect -1129 891 -1123 925
rect -1089 891 -1083 925
rect -1129 853 -1083 891
rect -1129 819 -1123 853
rect -1089 819 -1083 853
rect -1129 772 -1083 819
rect -971 925 -925 972
rect -971 891 -965 925
rect -931 891 -925 925
rect -971 853 -925 891
rect -971 819 -965 853
rect -931 819 -925 853
rect -971 772 -925 819
rect -813 925 -767 972
rect -813 891 -807 925
rect -773 891 -767 925
rect -813 853 -767 891
rect -813 819 -807 853
rect -773 819 -767 853
rect -813 772 -767 819
rect -655 925 -609 972
rect -655 891 -649 925
rect -615 891 -609 925
rect -655 853 -609 891
rect -655 819 -649 853
rect -615 819 -609 853
rect -655 772 -609 819
rect -497 925 -451 972
rect -497 891 -491 925
rect -457 891 -451 925
rect -497 853 -451 891
rect -497 819 -491 853
rect -457 819 -451 853
rect -497 772 -451 819
rect -339 925 -293 972
rect -339 891 -333 925
rect -299 891 -293 925
rect -339 853 -293 891
rect -339 819 -333 853
rect -299 819 -293 853
rect -339 772 -293 819
rect -181 925 -135 972
rect -181 891 -175 925
rect -141 891 -135 925
rect -181 853 -135 891
rect -181 819 -175 853
rect -141 819 -135 853
rect -181 772 -135 819
rect -23 925 23 972
rect -23 891 -17 925
rect 17 891 23 925
rect -23 853 23 891
rect -23 819 -17 853
rect 17 819 23 853
rect -23 772 23 819
rect 135 925 181 972
rect 135 891 141 925
rect 175 891 181 925
rect 135 853 181 891
rect 135 819 141 853
rect 175 819 181 853
rect 135 772 181 819
rect 293 925 339 972
rect 293 891 299 925
rect 333 891 339 925
rect 293 853 339 891
rect 293 819 299 853
rect 333 819 339 853
rect 293 772 339 819
rect 451 925 497 972
rect 451 891 457 925
rect 491 891 497 925
rect 451 853 497 891
rect 451 819 457 853
rect 491 819 497 853
rect 451 772 497 819
rect 609 925 655 972
rect 609 891 615 925
rect 649 891 655 925
rect 609 853 655 891
rect 609 819 615 853
rect 649 819 655 853
rect 609 772 655 819
rect 767 925 813 972
rect 767 891 773 925
rect 807 891 813 925
rect 767 853 813 891
rect 767 819 773 853
rect 807 819 813 853
rect 767 772 813 819
rect 925 925 971 972
rect 925 891 931 925
rect 965 891 971 925
rect 925 853 971 891
rect 925 819 931 853
rect 965 819 971 853
rect 925 772 971 819
rect 1083 925 1129 972
rect 1083 891 1089 925
rect 1123 891 1129 925
rect 1083 853 1129 891
rect 1083 819 1089 853
rect 1123 819 1129 853
rect 1083 772 1129 819
rect 1241 925 1287 972
rect 1241 891 1247 925
rect 1281 891 1287 925
rect 1241 853 1287 891
rect 1241 819 1247 853
rect 1281 819 1287 853
rect 1241 772 1287 819
rect 1399 925 1445 972
rect 1399 891 1405 925
rect 1439 891 1445 925
rect 1399 853 1445 891
rect 1399 819 1405 853
rect 1439 819 1445 853
rect 1399 772 1445 819
rect 1557 925 1603 972
rect 1557 891 1563 925
rect 1597 891 1603 925
rect 1557 853 1603 891
rect 1557 819 1563 853
rect 1597 819 1603 853
rect 1557 772 1603 819
rect 1715 925 1761 972
rect 1715 891 1721 925
rect 1755 891 1761 925
rect 1715 853 1761 891
rect 1715 819 1721 853
rect 1755 819 1761 853
rect 1715 772 1761 819
rect 1873 925 1919 972
rect 1873 891 1879 925
rect 1913 891 1919 925
rect 1873 853 1919 891
rect 1873 819 1879 853
rect 1913 819 1919 853
rect 1873 772 1919 819
rect 2031 925 2077 972
rect 2031 891 2037 925
rect 2071 891 2077 925
rect 2031 853 2077 891
rect 2031 819 2037 853
rect 2071 819 2077 853
rect 2031 772 2077 819
rect 2189 925 2235 972
rect 2189 891 2195 925
rect 2229 891 2235 925
rect 2189 853 2235 891
rect 2189 819 2195 853
rect 2229 819 2235 853
rect 2189 772 2235 819
rect 2347 925 2393 972
rect 2347 891 2353 925
rect 2387 891 2393 925
rect 2347 853 2393 891
rect 2347 819 2353 853
rect 2387 819 2393 853
rect 2347 772 2393 819
rect 2505 925 2551 972
rect 2505 891 2511 925
rect 2545 891 2551 925
rect 2505 853 2551 891
rect 2505 819 2511 853
rect 2545 819 2551 853
rect 2505 772 2551 819
rect 2663 925 2709 972
rect 2663 891 2669 925
rect 2703 891 2709 925
rect 2663 853 2709 891
rect 2663 819 2669 853
rect 2703 819 2709 853
rect 2663 772 2709 819
rect 2821 925 2867 972
rect 2821 891 2827 925
rect 2861 891 2867 925
rect 2821 853 2867 891
rect 2821 819 2827 853
rect 2861 819 2867 853
rect 2821 772 2867 819
rect 2979 925 3025 972
rect 2979 891 2985 925
rect 3019 891 3025 925
rect 2979 853 3025 891
rect 2979 819 2985 853
rect 3019 819 3025 853
rect 2979 772 3025 819
rect 3137 925 3183 972
rect 3137 891 3143 925
rect 3177 891 3183 925
rect 3137 853 3183 891
rect 3137 819 3143 853
rect 3177 819 3183 853
rect 3137 772 3183 819
rect -3127 725 -3035 731
rect -3127 691 -3098 725
rect -3064 691 -3035 725
rect -3127 685 -3035 691
rect -2969 725 -2877 731
rect -2969 691 -2940 725
rect -2906 691 -2877 725
rect -2969 685 -2877 691
rect -2811 725 -2719 731
rect -2811 691 -2782 725
rect -2748 691 -2719 725
rect -2811 685 -2719 691
rect -2653 725 -2561 731
rect -2653 691 -2624 725
rect -2590 691 -2561 725
rect -2653 685 -2561 691
rect -2495 725 -2403 731
rect -2495 691 -2466 725
rect -2432 691 -2403 725
rect -2495 685 -2403 691
rect -2337 725 -2245 731
rect -2337 691 -2308 725
rect -2274 691 -2245 725
rect -2337 685 -2245 691
rect -2179 725 -2087 731
rect -2179 691 -2150 725
rect -2116 691 -2087 725
rect -2179 685 -2087 691
rect -2021 725 -1929 731
rect -2021 691 -1992 725
rect -1958 691 -1929 725
rect -2021 685 -1929 691
rect -1863 725 -1771 731
rect -1863 691 -1834 725
rect -1800 691 -1771 725
rect -1863 685 -1771 691
rect -1705 725 -1613 731
rect -1705 691 -1676 725
rect -1642 691 -1613 725
rect -1705 685 -1613 691
rect -1547 725 -1455 731
rect -1547 691 -1518 725
rect -1484 691 -1455 725
rect -1547 685 -1455 691
rect -1389 725 -1297 731
rect -1389 691 -1360 725
rect -1326 691 -1297 725
rect -1389 685 -1297 691
rect -1231 725 -1139 731
rect -1231 691 -1202 725
rect -1168 691 -1139 725
rect -1231 685 -1139 691
rect -1073 725 -981 731
rect -1073 691 -1044 725
rect -1010 691 -981 725
rect -1073 685 -981 691
rect -915 725 -823 731
rect -915 691 -886 725
rect -852 691 -823 725
rect -915 685 -823 691
rect -757 725 -665 731
rect -757 691 -728 725
rect -694 691 -665 725
rect -757 685 -665 691
rect -599 725 -507 731
rect -599 691 -570 725
rect -536 691 -507 725
rect -599 685 -507 691
rect -441 725 -349 731
rect -441 691 -412 725
rect -378 691 -349 725
rect -441 685 -349 691
rect -283 725 -191 731
rect -283 691 -254 725
rect -220 691 -191 725
rect -283 685 -191 691
rect -125 725 -33 731
rect -125 691 -96 725
rect -62 691 -33 725
rect -125 685 -33 691
rect 33 725 125 731
rect 33 691 62 725
rect 96 691 125 725
rect 33 685 125 691
rect 191 725 283 731
rect 191 691 220 725
rect 254 691 283 725
rect 191 685 283 691
rect 349 725 441 731
rect 349 691 378 725
rect 412 691 441 725
rect 349 685 441 691
rect 507 725 599 731
rect 507 691 536 725
rect 570 691 599 725
rect 507 685 599 691
rect 665 725 757 731
rect 665 691 694 725
rect 728 691 757 725
rect 665 685 757 691
rect 823 725 915 731
rect 823 691 852 725
rect 886 691 915 725
rect 823 685 915 691
rect 981 725 1073 731
rect 981 691 1010 725
rect 1044 691 1073 725
rect 981 685 1073 691
rect 1139 725 1231 731
rect 1139 691 1168 725
rect 1202 691 1231 725
rect 1139 685 1231 691
rect 1297 725 1389 731
rect 1297 691 1326 725
rect 1360 691 1389 725
rect 1297 685 1389 691
rect 1455 725 1547 731
rect 1455 691 1484 725
rect 1518 691 1547 725
rect 1455 685 1547 691
rect 1613 725 1705 731
rect 1613 691 1642 725
rect 1676 691 1705 725
rect 1613 685 1705 691
rect 1771 725 1863 731
rect 1771 691 1800 725
rect 1834 691 1863 725
rect 1771 685 1863 691
rect 1929 725 2021 731
rect 1929 691 1958 725
rect 1992 691 2021 725
rect 1929 685 2021 691
rect 2087 725 2179 731
rect 2087 691 2116 725
rect 2150 691 2179 725
rect 2087 685 2179 691
rect 2245 725 2337 731
rect 2245 691 2274 725
rect 2308 691 2337 725
rect 2245 685 2337 691
rect 2403 725 2495 731
rect 2403 691 2432 725
rect 2466 691 2495 725
rect 2403 685 2495 691
rect 2561 725 2653 731
rect 2561 691 2590 725
rect 2624 691 2653 725
rect 2561 685 2653 691
rect 2719 725 2811 731
rect 2719 691 2748 725
rect 2782 691 2811 725
rect 2719 685 2811 691
rect 2877 725 2969 731
rect 2877 691 2906 725
rect 2940 691 2969 725
rect 2877 685 2969 691
rect 3035 725 3127 731
rect 3035 691 3064 725
rect 3098 691 3127 725
rect 3035 685 3127 691
rect -3127 617 -3035 623
rect -3127 583 -3098 617
rect -3064 583 -3035 617
rect -3127 577 -3035 583
rect -2969 617 -2877 623
rect -2969 583 -2940 617
rect -2906 583 -2877 617
rect -2969 577 -2877 583
rect -2811 617 -2719 623
rect -2811 583 -2782 617
rect -2748 583 -2719 617
rect -2811 577 -2719 583
rect -2653 617 -2561 623
rect -2653 583 -2624 617
rect -2590 583 -2561 617
rect -2653 577 -2561 583
rect -2495 617 -2403 623
rect -2495 583 -2466 617
rect -2432 583 -2403 617
rect -2495 577 -2403 583
rect -2337 617 -2245 623
rect -2337 583 -2308 617
rect -2274 583 -2245 617
rect -2337 577 -2245 583
rect -2179 617 -2087 623
rect -2179 583 -2150 617
rect -2116 583 -2087 617
rect -2179 577 -2087 583
rect -2021 617 -1929 623
rect -2021 583 -1992 617
rect -1958 583 -1929 617
rect -2021 577 -1929 583
rect -1863 617 -1771 623
rect -1863 583 -1834 617
rect -1800 583 -1771 617
rect -1863 577 -1771 583
rect -1705 617 -1613 623
rect -1705 583 -1676 617
rect -1642 583 -1613 617
rect -1705 577 -1613 583
rect -1547 617 -1455 623
rect -1547 583 -1518 617
rect -1484 583 -1455 617
rect -1547 577 -1455 583
rect -1389 617 -1297 623
rect -1389 583 -1360 617
rect -1326 583 -1297 617
rect -1389 577 -1297 583
rect -1231 617 -1139 623
rect -1231 583 -1202 617
rect -1168 583 -1139 617
rect -1231 577 -1139 583
rect -1073 617 -981 623
rect -1073 583 -1044 617
rect -1010 583 -981 617
rect -1073 577 -981 583
rect -915 617 -823 623
rect -915 583 -886 617
rect -852 583 -823 617
rect -915 577 -823 583
rect -757 617 -665 623
rect -757 583 -728 617
rect -694 583 -665 617
rect -757 577 -665 583
rect -599 617 -507 623
rect -599 583 -570 617
rect -536 583 -507 617
rect -599 577 -507 583
rect -441 617 -349 623
rect -441 583 -412 617
rect -378 583 -349 617
rect -441 577 -349 583
rect -283 617 -191 623
rect -283 583 -254 617
rect -220 583 -191 617
rect -283 577 -191 583
rect -125 617 -33 623
rect -125 583 -96 617
rect -62 583 -33 617
rect -125 577 -33 583
rect 33 617 125 623
rect 33 583 62 617
rect 96 583 125 617
rect 33 577 125 583
rect 191 617 283 623
rect 191 583 220 617
rect 254 583 283 617
rect 191 577 283 583
rect 349 617 441 623
rect 349 583 378 617
rect 412 583 441 617
rect 349 577 441 583
rect 507 617 599 623
rect 507 583 536 617
rect 570 583 599 617
rect 507 577 599 583
rect 665 617 757 623
rect 665 583 694 617
rect 728 583 757 617
rect 665 577 757 583
rect 823 617 915 623
rect 823 583 852 617
rect 886 583 915 617
rect 823 577 915 583
rect 981 617 1073 623
rect 981 583 1010 617
rect 1044 583 1073 617
rect 981 577 1073 583
rect 1139 617 1231 623
rect 1139 583 1168 617
rect 1202 583 1231 617
rect 1139 577 1231 583
rect 1297 617 1389 623
rect 1297 583 1326 617
rect 1360 583 1389 617
rect 1297 577 1389 583
rect 1455 617 1547 623
rect 1455 583 1484 617
rect 1518 583 1547 617
rect 1455 577 1547 583
rect 1613 617 1705 623
rect 1613 583 1642 617
rect 1676 583 1705 617
rect 1613 577 1705 583
rect 1771 617 1863 623
rect 1771 583 1800 617
rect 1834 583 1863 617
rect 1771 577 1863 583
rect 1929 617 2021 623
rect 1929 583 1958 617
rect 1992 583 2021 617
rect 1929 577 2021 583
rect 2087 617 2179 623
rect 2087 583 2116 617
rect 2150 583 2179 617
rect 2087 577 2179 583
rect 2245 617 2337 623
rect 2245 583 2274 617
rect 2308 583 2337 617
rect 2245 577 2337 583
rect 2403 617 2495 623
rect 2403 583 2432 617
rect 2466 583 2495 617
rect 2403 577 2495 583
rect 2561 617 2653 623
rect 2561 583 2590 617
rect 2624 583 2653 617
rect 2561 577 2653 583
rect 2719 617 2811 623
rect 2719 583 2748 617
rect 2782 583 2811 617
rect 2719 577 2811 583
rect 2877 617 2969 623
rect 2877 583 2906 617
rect 2940 583 2969 617
rect 2877 577 2969 583
rect 3035 617 3127 623
rect 3035 583 3064 617
rect 3098 583 3127 617
rect 3035 577 3127 583
rect -3183 489 -3137 536
rect -3183 455 -3177 489
rect -3143 455 -3137 489
rect -3183 417 -3137 455
rect -3183 383 -3177 417
rect -3143 383 -3137 417
rect -3183 336 -3137 383
rect -3025 489 -2979 536
rect -3025 455 -3019 489
rect -2985 455 -2979 489
rect -3025 417 -2979 455
rect -3025 383 -3019 417
rect -2985 383 -2979 417
rect -3025 336 -2979 383
rect -2867 489 -2821 536
rect -2867 455 -2861 489
rect -2827 455 -2821 489
rect -2867 417 -2821 455
rect -2867 383 -2861 417
rect -2827 383 -2821 417
rect -2867 336 -2821 383
rect -2709 489 -2663 536
rect -2709 455 -2703 489
rect -2669 455 -2663 489
rect -2709 417 -2663 455
rect -2709 383 -2703 417
rect -2669 383 -2663 417
rect -2709 336 -2663 383
rect -2551 489 -2505 536
rect -2551 455 -2545 489
rect -2511 455 -2505 489
rect -2551 417 -2505 455
rect -2551 383 -2545 417
rect -2511 383 -2505 417
rect -2551 336 -2505 383
rect -2393 489 -2347 536
rect -2393 455 -2387 489
rect -2353 455 -2347 489
rect -2393 417 -2347 455
rect -2393 383 -2387 417
rect -2353 383 -2347 417
rect -2393 336 -2347 383
rect -2235 489 -2189 536
rect -2235 455 -2229 489
rect -2195 455 -2189 489
rect -2235 417 -2189 455
rect -2235 383 -2229 417
rect -2195 383 -2189 417
rect -2235 336 -2189 383
rect -2077 489 -2031 536
rect -2077 455 -2071 489
rect -2037 455 -2031 489
rect -2077 417 -2031 455
rect -2077 383 -2071 417
rect -2037 383 -2031 417
rect -2077 336 -2031 383
rect -1919 489 -1873 536
rect -1919 455 -1913 489
rect -1879 455 -1873 489
rect -1919 417 -1873 455
rect -1919 383 -1913 417
rect -1879 383 -1873 417
rect -1919 336 -1873 383
rect -1761 489 -1715 536
rect -1761 455 -1755 489
rect -1721 455 -1715 489
rect -1761 417 -1715 455
rect -1761 383 -1755 417
rect -1721 383 -1715 417
rect -1761 336 -1715 383
rect -1603 489 -1557 536
rect -1603 455 -1597 489
rect -1563 455 -1557 489
rect -1603 417 -1557 455
rect -1603 383 -1597 417
rect -1563 383 -1557 417
rect -1603 336 -1557 383
rect -1445 489 -1399 536
rect -1445 455 -1439 489
rect -1405 455 -1399 489
rect -1445 417 -1399 455
rect -1445 383 -1439 417
rect -1405 383 -1399 417
rect -1445 336 -1399 383
rect -1287 489 -1241 536
rect -1287 455 -1281 489
rect -1247 455 -1241 489
rect -1287 417 -1241 455
rect -1287 383 -1281 417
rect -1247 383 -1241 417
rect -1287 336 -1241 383
rect -1129 489 -1083 536
rect -1129 455 -1123 489
rect -1089 455 -1083 489
rect -1129 417 -1083 455
rect -1129 383 -1123 417
rect -1089 383 -1083 417
rect -1129 336 -1083 383
rect -971 489 -925 536
rect -971 455 -965 489
rect -931 455 -925 489
rect -971 417 -925 455
rect -971 383 -965 417
rect -931 383 -925 417
rect -971 336 -925 383
rect -813 489 -767 536
rect -813 455 -807 489
rect -773 455 -767 489
rect -813 417 -767 455
rect -813 383 -807 417
rect -773 383 -767 417
rect -813 336 -767 383
rect -655 489 -609 536
rect -655 455 -649 489
rect -615 455 -609 489
rect -655 417 -609 455
rect -655 383 -649 417
rect -615 383 -609 417
rect -655 336 -609 383
rect -497 489 -451 536
rect -497 455 -491 489
rect -457 455 -451 489
rect -497 417 -451 455
rect -497 383 -491 417
rect -457 383 -451 417
rect -497 336 -451 383
rect -339 489 -293 536
rect -339 455 -333 489
rect -299 455 -293 489
rect -339 417 -293 455
rect -339 383 -333 417
rect -299 383 -293 417
rect -339 336 -293 383
rect -181 489 -135 536
rect -181 455 -175 489
rect -141 455 -135 489
rect -181 417 -135 455
rect -181 383 -175 417
rect -141 383 -135 417
rect -181 336 -135 383
rect -23 489 23 536
rect -23 455 -17 489
rect 17 455 23 489
rect -23 417 23 455
rect -23 383 -17 417
rect 17 383 23 417
rect -23 336 23 383
rect 135 489 181 536
rect 135 455 141 489
rect 175 455 181 489
rect 135 417 181 455
rect 135 383 141 417
rect 175 383 181 417
rect 135 336 181 383
rect 293 489 339 536
rect 293 455 299 489
rect 333 455 339 489
rect 293 417 339 455
rect 293 383 299 417
rect 333 383 339 417
rect 293 336 339 383
rect 451 489 497 536
rect 451 455 457 489
rect 491 455 497 489
rect 451 417 497 455
rect 451 383 457 417
rect 491 383 497 417
rect 451 336 497 383
rect 609 489 655 536
rect 609 455 615 489
rect 649 455 655 489
rect 609 417 655 455
rect 609 383 615 417
rect 649 383 655 417
rect 609 336 655 383
rect 767 489 813 536
rect 767 455 773 489
rect 807 455 813 489
rect 767 417 813 455
rect 767 383 773 417
rect 807 383 813 417
rect 767 336 813 383
rect 925 489 971 536
rect 925 455 931 489
rect 965 455 971 489
rect 925 417 971 455
rect 925 383 931 417
rect 965 383 971 417
rect 925 336 971 383
rect 1083 489 1129 536
rect 1083 455 1089 489
rect 1123 455 1129 489
rect 1083 417 1129 455
rect 1083 383 1089 417
rect 1123 383 1129 417
rect 1083 336 1129 383
rect 1241 489 1287 536
rect 1241 455 1247 489
rect 1281 455 1287 489
rect 1241 417 1287 455
rect 1241 383 1247 417
rect 1281 383 1287 417
rect 1241 336 1287 383
rect 1399 489 1445 536
rect 1399 455 1405 489
rect 1439 455 1445 489
rect 1399 417 1445 455
rect 1399 383 1405 417
rect 1439 383 1445 417
rect 1399 336 1445 383
rect 1557 489 1603 536
rect 1557 455 1563 489
rect 1597 455 1603 489
rect 1557 417 1603 455
rect 1557 383 1563 417
rect 1597 383 1603 417
rect 1557 336 1603 383
rect 1715 489 1761 536
rect 1715 455 1721 489
rect 1755 455 1761 489
rect 1715 417 1761 455
rect 1715 383 1721 417
rect 1755 383 1761 417
rect 1715 336 1761 383
rect 1873 489 1919 536
rect 1873 455 1879 489
rect 1913 455 1919 489
rect 1873 417 1919 455
rect 1873 383 1879 417
rect 1913 383 1919 417
rect 1873 336 1919 383
rect 2031 489 2077 536
rect 2031 455 2037 489
rect 2071 455 2077 489
rect 2031 417 2077 455
rect 2031 383 2037 417
rect 2071 383 2077 417
rect 2031 336 2077 383
rect 2189 489 2235 536
rect 2189 455 2195 489
rect 2229 455 2235 489
rect 2189 417 2235 455
rect 2189 383 2195 417
rect 2229 383 2235 417
rect 2189 336 2235 383
rect 2347 489 2393 536
rect 2347 455 2353 489
rect 2387 455 2393 489
rect 2347 417 2393 455
rect 2347 383 2353 417
rect 2387 383 2393 417
rect 2347 336 2393 383
rect 2505 489 2551 536
rect 2505 455 2511 489
rect 2545 455 2551 489
rect 2505 417 2551 455
rect 2505 383 2511 417
rect 2545 383 2551 417
rect 2505 336 2551 383
rect 2663 489 2709 536
rect 2663 455 2669 489
rect 2703 455 2709 489
rect 2663 417 2709 455
rect 2663 383 2669 417
rect 2703 383 2709 417
rect 2663 336 2709 383
rect 2821 489 2867 536
rect 2821 455 2827 489
rect 2861 455 2867 489
rect 2821 417 2867 455
rect 2821 383 2827 417
rect 2861 383 2867 417
rect 2821 336 2867 383
rect 2979 489 3025 536
rect 2979 455 2985 489
rect 3019 455 3025 489
rect 2979 417 3025 455
rect 2979 383 2985 417
rect 3019 383 3025 417
rect 2979 336 3025 383
rect 3137 489 3183 536
rect 3137 455 3143 489
rect 3177 455 3183 489
rect 3137 417 3183 455
rect 3137 383 3143 417
rect 3177 383 3183 417
rect 3137 336 3183 383
rect -3127 289 -3035 295
rect -3127 255 -3098 289
rect -3064 255 -3035 289
rect -3127 249 -3035 255
rect -2969 289 -2877 295
rect -2969 255 -2940 289
rect -2906 255 -2877 289
rect -2969 249 -2877 255
rect -2811 289 -2719 295
rect -2811 255 -2782 289
rect -2748 255 -2719 289
rect -2811 249 -2719 255
rect -2653 289 -2561 295
rect -2653 255 -2624 289
rect -2590 255 -2561 289
rect -2653 249 -2561 255
rect -2495 289 -2403 295
rect -2495 255 -2466 289
rect -2432 255 -2403 289
rect -2495 249 -2403 255
rect -2337 289 -2245 295
rect -2337 255 -2308 289
rect -2274 255 -2245 289
rect -2337 249 -2245 255
rect -2179 289 -2087 295
rect -2179 255 -2150 289
rect -2116 255 -2087 289
rect -2179 249 -2087 255
rect -2021 289 -1929 295
rect -2021 255 -1992 289
rect -1958 255 -1929 289
rect -2021 249 -1929 255
rect -1863 289 -1771 295
rect -1863 255 -1834 289
rect -1800 255 -1771 289
rect -1863 249 -1771 255
rect -1705 289 -1613 295
rect -1705 255 -1676 289
rect -1642 255 -1613 289
rect -1705 249 -1613 255
rect -1547 289 -1455 295
rect -1547 255 -1518 289
rect -1484 255 -1455 289
rect -1547 249 -1455 255
rect -1389 289 -1297 295
rect -1389 255 -1360 289
rect -1326 255 -1297 289
rect -1389 249 -1297 255
rect -1231 289 -1139 295
rect -1231 255 -1202 289
rect -1168 255 -1139 289
rect -1231 249 -1139 255
rect -1073 289 -981 295
rect -1073 255 -1044 289
rect -1010 255 -981 289
rect -1073 249 -981 255
rect -915 289 -823 295
rect -915 255 -886 289
rect -852 255 -823 289
rect -915 249 -823 255
rect -757 289 -665 295
rect -757 255 -728 289
rect -694 255 -665 289
rect -757 249 -665 255
rect -599 289 -507 295
rect -599 255 -570 289
rect -536 255 -507 289
rect -599 249 -507 255
rect -441 289 -349 295
rect -441 255 -412 289
rect -378 255 -349 289
rect -441 249 -349 255
rect -283 289 -191 295
rect -283 255 -254 289
rect -220 255 -191 289
rect -283 249 -191 255
rect -125 289 -33 295
rect -125 255 -96 289
rect -62 255 -33 289
rect -125 249 -33 255
rect 33 289 125 295
rect 33 255 62 289
rect 96 255 125 289
rect 33 249 125 255
rect 191 289 283 295
rect 191 255 220 289
rect 254 255 283 289
rect 191 249 283 255
rect 349 289 441 295
rect 349 255 378 289
rect 412 255 441 289
rect 349 249 441 255
rect 507 289 599 295
rect 507 255 536 289
rect 570 255 599 289
rect 507 249 599 255
rect 665 289 757 295
rect 665 255 694 289
rect 728 255 757 289
rect 665 249 757 255
rect 823 289 915 295
rect 823 255 852 289
rect 886 255 915 289
rect 823 249 915 255
rect 981 289 1073 295
rect 981 255 1010 289
rect 1044 255 1073 289
rect 981 249 1073 255
rect 1139 289 1231 295
rect 1139 255 1168 289
rect 1202 255 1231 289
rect 1139 249 1231 255
rect 1297 289 1389 295
rect 1297 255 1326 289
rect 1360 255 1389 289
rect 1297 249 1389 255
rect 1455 289 1547 295
rect 1455 255 1484 289
rect 1518 255 1547 289
rect 1455 249 1547 255
rect 1613 289 1705 295
rect 1613 255 1642 289
rect 1676 255 1705 289
rect 1613 249 1705 255
rect 1771 289 1863 295
rect 1771 255 1800 289
rect 1834 255 1863 289
rect 1771 249 1863 255
rect 1929 289 2021 295
rect 1929 255 1958 289
rect 1992 255 2021 289
rect 1929 249 2021 255
rect 2087 289 2179 295
rect 2087 255 2116 289
rect 2150 255 2179 289
rect 2087 249 2179 255
rect 2245 289 2337 295
rect 2245 255 2274 289
rect 2308 255 2337 289
rect 2245 249 2337 255
rect 2403 289 2495 295
rect 2403 255 2432 289
rect 2466 255 2495 289
rect 2403 249 2495 255
rect 2561 289 2653 295
rect 2561 255 2590 289
rect 2624 255 2653 289
rect 2561 249 2653 255
rect 2719 289 2811 295
rect 2719 255 2748 289
rect 2782 255 2811 289
rect 2719 249 2811 255
rect 2877 289 2969 295
rect 2877 255 2906 289
rect 2940 255 2969 289
rect 2877 249 2969 255
rect 3035 289 3127 295
rect 3035 255 3064 289
rect 3098 255 3127 289
rect 3035 249 3127 255
rect -3127 181 -3035 187
rect -3127 147 -3098 181
rect -3064 147 -3035 181
rect -3127 141 -3035 147
rect -2969 181 -2877 187
rect -2969 147 -2940 181
rect -2906 147 -2877 181
rect -2969 141 -2877 147
rect -2811 181 -2719 187
rect -2811 147 -2782 181
rect -2748 147 -2719 181
rect -2811 141 -2719 147
rect -2653 181 -2561 187
rect -2653 147 -2624 181
rect -2590 147 -2561 181
rect -2653 141 -2561 147
rect -2495 181 -2403 187
rect -2495 147 -2466 181
rect -2432 147 -2403 181
rect -2495 141 -2403 147
rect -2337 181 -2245 187
rect -2337 147 -2308 181
rect -2274 147 -2245 181
rect -2337 141 -2245 147
rect -2179 181 -2087 187
rect -2179 147 -2150 181
rect -2116 147 -2087 181
rect -2179 141 -2087 147
rect -2021 181 -1929 187
rect -2021 147 -1992 181
rect -1958 147 -1929 181
rect -2021 141 -1929 147
rect -1863 181 -1771 187
rect -1863 147 -1834 181
rect -1800 147 -1771 181
rect -1863 141 -1771 147
rect -1705 181 -1613 187
rect -1705 147 -1676 181
rect -1642 147 -1613 181
rect -1705 141 -1613 147
rect -1547 181 -1455 187
rect -1547 147 -1518 181
rect -1484 147 -1455 181
rect -1547 141 -1455 147
rect -1389 181 -1297 187
rect -1389 147 -1360 181
rect -1326 147 -1297 181
rect -1389 141 -1297 147
rect -1231 181 -1139 187
rect -1231 147 -1202 181
rect -1168 147 -1139 181
rect -1231 141 -1139 147
rect -1073 181 -981 187
rect -1073 147 -1044 181
rect -1010 147 -981 181
rect -1073 141 -981 147
rect -915 181 -823 187
rect -915 147 -886 181
rect -852 147 -823 181
rect -915 141 -823 147
rect -757 181 -665 187
rect -757 147 -728 181
rect -694 147 -665 181
rect -757 141 -665 147
rect -599 181 -507 187
rect -599 147 -570 181
rect -536 147 -507 181
rect -599 141 -507 147
rect -441 181 -349 187
rect -441 147 -412 181
rect -378 147 -349 181
rect -441 141 -349 147
rect -283 181 -191 187
rect -283 147 -254 181
rect -220 147 -191 181
rect -283 141 -191 147
rect -125 181 -33 187
rect -125 147 -96 181
rect -62 147 -33 181
rect -125 141 -33 147
rect 33 181 125 187
rect 33 147 62 181
rect 96 147 125 181
rect 33 141 125 147
rect 191 181 283 187
rect 191 147 220 181
rect 254 147 283 181
rect 191 141 283 147
rect 349 181 441 187
rect 349 147 378 181
rect 412 147 441 181
rect 349 141 441 147
rect 507 181 599 187
rect 507 147 536 181
rect 570 147 599 181
rect 507 141 599 147
rect 665 181 757 187
rect 665 147 694 181
rect 728 147 757 181
rect 665 141 757 147
rect 823 181 915 187
rect 823 147 852 181
rect 886 147 915 181
rect 823 141 915 147
rect 981 181 1073 187
rect 981 147 1010 181
rect 1044 147 1073 181
rect 981 141 1073 147
rect 1139 181 1231 187
rect 1139 147 1168 181
rect 1202 147 1231 181
rect 1139 141 1231 147
rect 1297 181 1389 187
rect 1297 147 1326 181
rect 1360 147 1389 181
rect 1297 141 1389 147
rect 1455 181 1547 187
rect 1455 147 1484 181
rect 1518 147 1547 181
rect 1455 141 1547 147
rect 1613 181 1705 187
rect 1613 147 1642 181
rect 1676 147 1705 181
rect 1613 141 1705 147
rect 1771 181 1863 187
rect 1771 147 1800 181
rect 1834 147 1863 181
rect 1771 141 1863 147
rect 1929 181 2021 187
rect 1929 147 1958 181
rect 1992 147 2021 181
rect 1929 141 2021 147
rect 2087 181 2179 187
rect 2087 147 2116 181
rect 2150 147 2179 181
rect 2087 141 2179 147
rect 2245 181 2337 187
rect 2245 147 2274 181
rect 2308 147 2337 181
rect 2245 141 2337 147
rect 2403 181 2495 187
rect 2403 147 2432 181
rect 2466 147 2495 181
rect 2403 141 2495 147
rect 2561 181 2653 187
rect 2561 147 2590 181
rect 2624 147 2653 181
rect 2561 141 2653 147
rect 2719 181 2811 187
rect 2719 147 2748 181
rect 2782 147 2811 181
rect 2719 141 2811 147
rect 2877 181 2969 187
rect 2877 147 2906 181
rect 2940 147 2969 181
rect 2877 141 2969 147
rect 3035 181 3127 187
rect 3035 147 3064 181
rect 3098 147 3127 181
rect 3035 141 3127 147
rect -3183 53 -3137 100
rect -3183 19 -3177 53
rect -3143 19 -3137 53
rect -3183 -19 -3137 19
rect -3183 -53 -3177 -19
rect -3143 -53 -3137 -19
rect -3183 -100 -3137 -53
rect -3025 53 -2979 100
rect -3025 19 -3019 53
rect -2985 19 -2979 53
rect -3025 -19 -2979 19
rect -3025 -53 -3019 -19
rect -2985 -53 -2979 -19
rect -3025 -100 -2979 -53
rect -2867 53 -2821 100
rect -2867 19 -2861 53
rect -2827 19 -2821 53
rect -2867 -19 -2821 19
rect -2867 -53 -2861 -19
rect -2827 -53 -2821 -19
rect -2867 -100 -2821 -53
rect -2709 53 -2663 100
rect -2709 19 -2703 53
rect -2669 19 -2663 53
rect -2709 -19 -2663 19
rect -2709 -53 -2703 -19
rect -2669 -53 -2663 -19
rect -2709 -100 -2663 -53
rect -2551 53 -2505 100
rect -2551 19 -2545 53
rect -2511 19 -2505 53
rect -2551 -19 -2505 19
rect -2551 -53 -2545 -19
rect -2511 -53 -2505 -19
rect -2551 -100 -2505 -53
rect -2393 53 -2347 100
rect -2393 19 -2387 53
rect -2353 19 -2347 53
rect -2393 -19 -2347 19
rect -2393 -53 -2387 -19
rect -2353 -53 -2347 -19
rect -2393 -100 -2347 -53
rect -2235 53 -2189 100
rect -2235 19 -2229 53
rect -2195 19 -2189 53
rect -2235 -19 -2189 19
rect -2235 -53 -2229 -19
rect -2195 -53 -2189 -19
rect -2235 -100 -2189 -53
rect -2077 53 -2031 100
rect -2077 19 -2071 53
rect -2037 19 -2031 53
rect -2077 -19 -2031 19
rect -2077 -53 -2071 -19
rect -2037 -53 -2031 -19
rect -2077 -100 -2031 -53
rect -1919 53 -1873 100
rect -1919 19 -1913 53
rect -1879 19 -1873 53
rect -1919 -19 -1873 19
rect -1919 -53 -1913 -19
rect -1879 -53 -1873 -19
rect -1919 -100 -1873 -53
rect -1761 53 -1715 100
rect -1761 19 -1755 53
rect -1721 19 -1715 53
rect -1761 -19 -1715 19
rect -1761 -53 -1755 -19
rect -1721 -53 -1715 -19
rect -1761 -100 -1715 -53
rect -1603 53 -1557 100
rect -1603 19 -1597 53
rect -1563 19 -1557 53
rect -1603 -19 -1557 19
rect -1603 -53 -1597 -19
rect -1563 -53 -1557 -19
rect -1603 -100 -1557 -53
rect -1445 53 -1399 100
rect -1445 19 -1439 53
rect -1405 19 -1399 53
rect -1445 -19 -1399 19
rect -1445 -53 -1439 -19
rect -1405 -53 -1399 -19
rect -1445 -100 -1399 -53
rect -1287 53 -1241 100
rect -1287 19 -1281 53
rect -1247 19 -1241 53
rect -1287 -19 -1241 19
rect -1287 -53 -1281 -19
rect -1247 -53 -1241 -19
rect -1287 -100 -1241 -53
rect -1129 53 -1083 100
rect -1129 19 -1123 53
rect -1089 19 -1083 53
rect -1129 -19 -1083 19
rect -1129 -53 -1123 -19
rect -1089 -53 -1083 -19
rect -1129 -100 -1083 -53
rect -971 53 -925 100
rect -971 19 -965 53
rect -931 19 -925 53
rect -971 -19 -925 19
rect -971 -53 -965 -19
rect -931 -53 -925 -19
rect -971 -100 -925 -53
rect -813 53 -767 100
rect -813 19 -807 53
rect -773 19 -767 53
rect -813 -19 -767 19
rect -813 -53 -807 -19
rect -773 -53 -767 -19
rect -813 -100 -767 -53
rect -655 53 -609 100
rect -655 19 -649 53
rect -615 19 -609 53
rect -655 -19 -609 19
rect -655 -53 -649 -19
rect -615 -53 -609 -19
rect -655 -100 -609 -53
rect -497 53 -451 100
rect -497 19 -491 53
rect -457 19 -451 53
rect -497 -19 -451 19
rect -497 -53 -491 -19
rect -457 -53 -451 -19
rect -497 -100 -451 -53
rect -339 53 -293 100
rect -339 19 -333 53
rect -299 19 -293 53
rect -339 -19 -293 19
rect -339 -53 -333 -19
rect -299 -53 -293 -19
rect -339 -100 -293 -53
rect -181 53 -135 100
rect -181 19 -175 53
rect -141 19 -135 53
rect -181 -19 -135 19
rect -181 -53 -175 -19
rect -141 -53 -135 -19
rect -181 -100 -135 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 135 53 181 100
rect 135 19 141 53
rect 175 19 181 53
rect 135 -19 181 19
rect 135 -53 141 -19
rect 175 -53 181 -19
rect 135 -100 181 -53
rect 293 53 339 100
rect 293 19 299 53
rect 333 19 339 53
rect 293 -19 339 19
rect 293 -53 299 -19
rect 333 -53 339 -19
rect 293 -100 339 -53
rect 451 53 497 100
rect 451 19 457 53
rect 491 19 497 53
rect 451 -19 497 19
rect 451 -53 457 -19
rect 491 -53 497 -19
rect 451 -100 497 -53
rect 609 53 655 100
rect 609 19 615 53
rect 649 19 655 53
rect 609 -19 655 19
rect 609 -53 615 -19
rect 649 -53 655 -19
rect 609 -100 655 -53
rect 767 53 813 100
rect 767 19 773 53
rect 807 19 813 53
rect 767 -19 813 19
rect 767 -53 773 -19
rect 807 -53 813 -19
rect 767 -100 813 -53
rect 925 53 971 100
rect 925 19 931 53
rect 965 19 971 53
rect 925 -19 971 19
rect 925 -53 931 -19
rect 965 -53 971 -19
rect 925 -100 971 -53
rect 1083 53 1129 100
rect 1083 19 1089 53
rect 1123 19 1129 53
rect 1083 -19 1129 19
rect 1083 -53 1089 -19
rect 1123 -53 1129 -19
rect 1083 -100 1129 -53
rect 1241 53 1287 100
rect 1241 19 1247 53
rect 1281 19 1287 53
rect 1241 -19 1287 19
rect 1241 -53 1247 -19
rect 1281 -53 1287 -19
rect 1241 -100 1287 -53
rect 1399 53 1445 100
rect 1399 19 1405 53
rect 1439 19 1445 53
rect 1399 -19 1445 19
rect 1399 -53 1405 -19
rect 1439 -53 1445 -19
rect 1399 -100 1445 -53
rect 1557 53 1603 100
rect 1557 19 1563 53
rect 1597 19 1603 53
rect 1557 -19 1603 19
rect 1557 -53 1563 -19
rect 1597 -53 1603 -19
rect 1557 -100 1603 -53
rect 1715 53 1761 100
rect 1715 19 1721 53
rect 1755 19 1761 53
rect 1715 -19 1761 19
rect 1715 -53 1721 -19
rect 1755 -53 1761 -19
rect 1715 -100 1761 -53
rect 1873 53 1919 100
rect 1873 19 1879 53
rect 1913 19 1919 53
rect 1873 -19 1919 19
rect 1873 -53 1879 -19
rect 1913 -53 1919 -19
rect 1873 -100 1919 -53
rect 2031 53 2077 100
rect 2031 19 2037 53
rect 2071 19 2077 53
rect 2031 -19 2077 19
rect 2031 -53 2037 -19
rect 2071 -53 2077 -19
rect 2031 -100 2077 -53
rect 2189 53 2235 100
rect 2189 19 2195 53
rect 2229 19 2235 53
rect 2189 -19 2235 19
rect 2189 -53 2195 -19
rect 2229 -53 2235 -19
rect 2189 -100 2235 -53
rect 2347 53 2393 100
rect 2347 19 2353 53
rect 2387 19 2393 53
rect 2347 -19 2393 19
rect 2347 -53 2353 -19
rect 2387 -53 2393 -19
rect 2347 -100 2393 -53
rect 2505 53 2551 100
rect 2505 19 2511 53
rect 2545 19 2551 53
rect 2505 -19 2551 19
rect 2505 -53 2511 -19
rect 2545 -53 2551 -19
rect 2505 -100 2551 -53
rect 2663 53 2709 100
rect 2663 19 2669 53
rect 2703 19 2709 53
rect 2663 -19 2709 19
rect 2663 -53 2669 -19
rect 2703 -53 2709 -19
rect 2663 -100 2709 -53
rect 2821 53 2867 100
rect 2821 19 2827 53
rect 2861 19 2867 53
rect 2821 -19 2867 19
rect 2821 -53 2827 -19
rect 2861 -53 2867 -19
rect 2821 -100 2867 -53
rect 2979 53 3025 100
rect 2979 19 2985 53
rect 3019 19 3025 53
rect 2979 -19 3025 19
rect 2979 -53 2985 -19
rect 3019 -53 3025 -19
rect 2979 -100 3025 -53
rect 3137 53 3183 100
rect 3137 19 3143 53
rect 3177 19 3183 53
rect 3137 -19 3183 19
rect 3137 -53 3143 -19
rect 3177 -53 3183 -19
rect 3137 -100 3183 -53
rect -3127 -147 -3035 -141
rect -3127 -181 -3098 -147
rect -3064 -181 -3035 -147
rect -3127 -187 -3035 -181
rect -2969 -147 -2877 -141
rect -2969 -181 -2940 -147
rect -2906 -181 -2877 -147
rect -2969 -187 -2877 -181
rect -2811 -147 -2719 -141
rect -2811 -181 -2782 -147
rect -2748 -181 -2719 -147
rect -2811 -187 -2719 -181
rect -2653 -147 -2561 -141
rect -2653 -181 -2624 -147
rect -2590 -181 -2561 -147
rect -2653 -187 -2561 -181
rect -2495 -147 -2403 -141
rect -2495 -181 -2466 -147
rect -2432 -181 -2403 -147
rect -2495 -187 -2403 -181
rect -2337 -147 -2245 -141
rect -2337 -181 -2308 -147
rect -2274 -181 -2245 -147
rect -2337 -187 -2245 -181
rect -2179 -147 -2087 -141
rect -2179 -181 -2150 -147
rect -2116 -181 -2087 -147
rect -2179 -187 -2087 -181
rect -2021 -147 -1929 -141
rect -2021 -181 -1992 -147
rect -1958 -181 -1929 -147
rect -2021 -187 -1929 -181
rect -1863 -147 -1771 -141
rect -1863 -181 -1834 -147
rect -1800 -181 -1771 -147
rect -1863 -187 -1771 -181
rect -1705 -147 -1613 -141
rect -1705 -181 -1676 -147
rect -1642 -181 -1613 -147
rect -1705 -187 -1613 -181
rect -1547 -147 -1455 -141
rect -1547 -181 -1518 -147
rect -1484 -181 -1455 -147
rect -1547 -187 -1455 -181
rect -1389 -147 -1297 -141
rect -1389 -181 -1360 -147
rect -1326 -181 -1297 -147
rect -1389 -187 -1297 -181
rect -1231 -147 -1139 -141
rect -1231 -181 -1202 -147
rect -1168 -181 -1139 -147
rect -1231 -187 -1139 -181
rect -1073 -147 -981 -141
rect -1073 -181 -1044 -147
rect -1010 -181 -981 -147
rect -1073 -187 -981 -181
rect -915 -147 -823 -141
rect -915 -181 -886 -147
rect -852 -181 -823 -147
rect -915 -187 -823 -181
rect -757 -147 -665 -141
rect -757 -181 -728 -147
rect -694 -181 -665 -147
rect -757 -187 -665 -181
rect -599 -147 -507 -141
rect -599 -181 -570 -147
rect -536 -181 -507 -147
rect -599 -187 -507 -181
rect -441 -147 -349 -141
rect -441 -181 -412 -147
rect -378 -181 -349 -147
rect -441 -187 -349 -181
rect -283 -147 -191 -141
rect -283 -181 -254 -147
rect -220 -181 -191 -147
rect -283 -187 -191 -181
rect -125 -147 -33 -141
rect -125 -181 -96 -147
rect -62 -181 -33 -147
rect -125 -187 -33 -181
rect 33 -147 125 -141
rect 33 -181 62 -147
rect 96 -181 125 -147
rect 33 -187 125 -181
rect 191 -147 283 -141
rect 191 -181 220 -147
rect 254 -181 283 -147
rect 191 -187 283 -181
rect 349 -147 441 -141
rect 349 -181 378 -147
rect 412 -181 441 -147
rect 349 -187 441 -181
rect 507 -147 599 -141
rect 507 -181 536 -147
rect 570 -181 599 -147
rect 507 -187 599 -181
rect 665 -147 757 -141
rect 665 -181 694 -147
rect 728 -181 757 -147
rect 665 -187 757 -181
rect 823 -147 915 -141
rect 823 -181 852 -147
rect 886 -181 915 -147
rect 823 -187 915 -181
rect 981 -147 1073 -141
rect 981 -181 1010 -147
rect 1044 -181 1073 -147
rect 981 -187 1073 -181
rect 1139 -147 1231 -141
rect 1139 -181 1168 -147
rect 1202 -181 1231 -147
rect 1139 -187 1231 -181
rect 1297 -147 1389 -141
rect 1297 -181 1326 -147
rect 1360 -181 1389 -147
rect 1297 -187 1389 -181
rect 1455 -147 1547 -141
rect 1455 -181 1484 -147
rect 1518 -181 1547 -147
rect 1455 -187 1547 -181
rect 1613 -147 1705 -141
rect 1613 -181 1642 -147
rect 1676 -181 1705 -147
rect 1613 -187 1705 -181
rect 1771 -147 1863 -141
rect 1771 -181 1800 -147
rect 1834 -181 1863 -147
rect 1771 -187 1863 -181
rect 1929 -147 2021 -141
rect 1929 -181 1958 -147
rect 1992 -181 2021 -147
rect 1929 -187 2021 -181
rect 2087 -147 2179 -141
rect 2087 -181 2116 -147
rect 2150 -181 2179 -147
rect 2087 -187 2179 -181
rect 2245 -147 2337 -141
rect 2245 -181 2274 -147
rect 2308 -181 2337 -147
rect 2245 -187 2337 -181
rect 2403 -147 2495 -141
rect 2403 -181 2432 -147
rect 2466 -181 2495 -147
rect 2403 -187 2495 -181
rect 2561 -147 2653 -141
rect 2561 -181 2590 -147
rect 2624 -181 2653 -147
rect 2561 -187 2653 -181
rect 2719 -147 2811 -141
rect 2719 -181 2748 -147
rect 2782 -181 2811 -147
rect 2719 -187 2811 -181
rect 2877 -147 2969 -141
rect 2877 -181 2906 -147
rect 2940 -181 2969 -147
rect 2877 -187 2969 -181
rect 3035 -147 3127 -141
rect 3035 -181 3064 -147
rect 3098 -181 3127 -147
rect 3035 -187 3127 -181
rect -3127 -255 -3035 -249
rect -3127 -289 -3098 -255
rect -3064 -289 -3035 -255
rect -3127 -295 -3035 -289
rect -2969 -255 -2877 -249
rect -2969 -289 -2940 -255
rect -2906 -289 -2877 -255
rect -2969 -295 -2877 -289
rect -2811 -255 -2719 -249
rect -2811 -289 -2782 -255
rect -2748 -289 -2719 -255
rect -2811 -295 -2719 -289
rect -2653 -255 -2561 -249
rect -2653 -289 -2624 -255
rect -2590 -289 -2561 -255
rect -2653 -295 -2561 -289
rect -2495 -255 -2403 -249
rect -2495 -289 -2466 -255
rect -2432 -289 -2403 -255
rect -2495 -295 -2403 -289
rect -2337 -255 -2245 -249
rect -2337 -289 -2308 -255
rect -2274 -289 -2245 -255
rect -2337 -295 -2245 -289
rect -2179 -255 -2087 -249
rect -2179 -289 -2150 -255
rect -2116 -289 -2087 -255
rect -2179 -295 -2087 -289
rect -2021 -255 -1929 -249
rect -2021 -289 -1992 -255
rect -1958 -289 -1929 -255
rect -2021 -295 -1929 -289
rect -1863 -255 -1771 -249
rect -1863 -289 -1834 -255
rect -1800 -289 -1771 -255
rect -1863 -295 -1771 -289
rect -1705 -255 -1613 -249
rect -1705 -289 -1676 -255
rect -1642 -289 -1613 -255
rect -1705 -295 -1613 -289
rect -1547 -255 -1455 -249
rect -1547 -289 -1518 -255
rect -1484 -289 -1455 -255
rect -1547 -295 -1455 -289
rect -1389 -255 -1297 -249
rect -1389 -289 -1360 -255
rect -1326 -289 -1297 -255
rect -1389 -295 -1297 -289
rect -1231 -255 -1139 -249
rect -1231 -289 -1202 -255
rect -1168 -289 -1139 -255
rect -1231 -295 -1139 -289
rect -1073 -255 -981 -249
rect -1073 -289 -1044 -255
rect -1010 -289 -981 -255
rect -1073 -295 -981 -289
rect -915 -255 -823 -249
rect -915 -289 -886 -255
rect -852 -289 -823 -255
rect -915 -295 -823 -289
rect -757 -255 -665 -249
rect -757 -289 -728 -255
rect -694 -289 -665 -255
rect -757 -295 -665 -289
rect -599 -255 -507 -249
rect -599 -289 -570 -255
rect -536 -289 -507 -255
rect -599 -295 -507 -289
rect -441 -255 -349 -249
rect -441 -289 -412 -255
rect -378 -289 -349 -255
rect -441 -295 -349 -289
rect -283 -255 -191 -249
rect -283 -289 -254 -255
rect -220 -289 -191 -255
rect -283 -295 -191 -289
rect -125 -255 -33 -249
rect -125 -289 -96 -255
rect -62 -289 -33 -255
rect -125 -295 -33 -289
rect 33 -255 125 -249
rect 33 -289 62 -255
rect 96 -289 125 -255
rect 33 -295 125 -289
rect 191 -255 283 -249
rect 191 -289 220 -255
rect 254 -289 283 -255
rect 191 -295 283 -289
rect 349 -255 441 -249
rect 349 -289 378 -255
rect 412 -289 441 -255
rect 349 -295 441 -289
rect 507 -255 599 -249
rect 507 -289 536 -255
rect 570 -289 599 -255
rect 507 -295 599 -289
rect 665 -255 757 -249
rect 665 -289 694 -255
rect 728 -289 757 -255
rect 665 -295 757 -289
rect 823 -255 915 -249
rect 823 -289 852 -255
rect 886 -289 915 -255
rect 823 -295 915 -289
rect 981 -255 1073 -249
rect 981 -289 1010 -255
rect 1044 -289 1073 -255
rect 981 -295 1073 -289
rect 1139 -255 1231 -249
rect 1139 -289 1168 -255
rect 1202 -289 1231 -255
rect 1139 -295 1231 -289
rect 1297 -255 1389 -249
rect 1297 -289 1326 -255
rect 1360 -289 1389 -255
rect 1297 -295 1389 -289
rect 1455 -255 1547 -249
rect 1455 -289 1484 -255
rect 1518 -289 1547 -255
rect 1455 -295 1547 -289
rect 1613 -255 1705 -249
rect 1613 -289 1642 -255
rect 1676 -289 1705 -255
rect 1613 -295 1705 -289
rect 1771 -255 1863 -249
rect 1771 -289 1800 -255
rect 1834 -289 1863 -255
rect 1771 -295 1863 -289
rect 1929 -255 2021 -249
rect 1929 -289 1958 -255
rect 1992 -289 2021 -255
rect 1929 -295 2021 -289
rect 2087 -255 2179 -249
rect 2087 -289 2116 -255
rect 2150 -289 2179 -255
rect 2087 -295 2179 -289
rect 2245 -255 2337 -249
rect 2245 -289 2274 -255
rect 2308 -289 2337 -255
rect 2245 -295 2337 -289
rect 2403 -255 2495 -249
rect 2403 -289 2432 -255
rect 2466 -289 2495 -255
rect 2403 -295 2495 -289
rect 2561 -255 2653 -249
rect 2561 -289 2590 -255
rect 2624 -289 2653 -255
rect 2561 -295 2653 -289
rect 2719 -255 2811 -249
rect 2719 -289 2748 -255
rect 2782 -289 2811 -255
rect 2719 -295 2811 -289
rect 2877 -255 2969 -249
rect 2877 -289 2906 -255
rect 2940 -289 2969 -255
rect 2877 -295 2969 -289
rect 3035 -255 3127 -249
rect 3035 -289 3064 -255
rect 3098 -289 3127 -255
rect 3035 -295 3127 -289
rect -3183 -383 -3137 -336
rect -3183 -417 -3177 -383
rect -3143 -417 -3137 -383
rect -3183 -455 -3137 -417
rect -3183 -489 -3177 -455
rect -3143 -489 -3137 -455
rect -3183 -536 -3137 -489
rect -3025 -383 -2979 -336
rect -3025 -417 -3019 -383
rect -2985 -417 -2979 -383
rect -3025 -455 -2979 -417
rect -3025 -489 -3019 -455
rect -2985 -489 -2979 -455
rect -3025 -536 -2979 -489
rect -2867 -383 -2821 -336
rect -2867 -417 -2861 -383
rect -2827 -417 -2821 -383
rect -2867 -455 -2821 -417
rect -2867 -489 -2861 -455
rect -2827 -489 -2821 -455
rect -2867 -536 -2821 -489
rect -2709 -383 -2663 -336
rect -2709 -417 -2703 -383
rect -2669 -417 -2663 -383
rect -2709 -455 -2663 -417
rect -2709 -489 -2703 -455
rect -2669 -489 -2663 -455
rect -2709 -536 -2663 -489
rect -2551 -383 -2505 -336
rect -2551 -417 -2545 -383
rect -2511 -417 -2505 -383
rect -2551 -455 -2505 -417
rect -2551 -489 -2545 -455
rect -2511 -489 -2505 -455
rect -2551 -536 -2505 -489
rect -2393 -383 -2347 -336
rect -2393 -417 -2387 -383
rect -2353 -417 -2347 -383
rect -2393 -455 -2347 -417
rect -2393 -489 -2387 -455
rect -2353 -489 -2347 -455
rect -2393 -536 -2347 -489
rect -2235 -383 -2189 -336
rect -2235 -417 -2229 -383
rect -2195 -417 -2189 -383
rect -2235 -455 -2189 -417
rect -2235 -489 -2229 -455
rect -2195 -489 -2189 -455
rect -2235 -536 -2189 -489
rect -2077 -383 -2031 -336
rect -2077 -417 -2071 -383
rect -2037 -417 -2031 -383
rect -2077 -455 -2031 -417
rect -2077 -489 -2071 -455
rect -2037 -489 -2031 -455
rect -2077 -536 -2031 -489
rect -1919 -383 -1873 -336
rect -1919 -417 -1913 -383
rect -1879 -417 -1873 -383
rect -1919 -455 -1873 -417
rect -1919 -489 -1913 -455
rect -1879 -489 -1873 -455
rect -1919 -536 -1873 -489
rect -1761 -383 -1715 -336
rect -1761 -417 -1755 -383
rect -1721 -417 -1715 -383
rect -1761 -455 -1715 -417
rect -1761 -489 -1755 -455
rect -1721 -489 -1715 -455
rect -1761 -536 -1715 -489
rect -1603 -383 -1557 -336
rect -1603 -417 -1597 -383
rect -1563 -417 -1557 -383
rect -1603 -455 -1557 -417
rect -1603 -489 -1597 -455
rect -1563 -489 -1557 -455
rect -1603 -536 -1557 -489
rect -1445 -383 -1399 -336
rect -1445 -417 -1439 -383
rect -1405 -417 -1399 -383
rect -1445 -455 -1399 -417
rect -1445 -489 -1439 -455
rect -1405 -489 -1399 -455
rect -1445 -536 -1399 -489
rect -1287 -383 -1241 -336
rect -1287 -417 -1281 -383
rect -1247 -417 -1241 -383
rect -1287 -455 -1241 -417
rect -1287 -489 -1281 -455
rect -1247 -489 -1241 -455
rect -1287 -536 -1241 -489
rect -1129 -383 -1083 -336
rect -1129 -417 -1123 -383
rect -1089 -417 -1083 -383
rect -1129 -455 -1083 -417
rect -1129 -489 -1123 -455
rect -1089 -489 -1083 -455
rect -1129 -536 -1083 -489
rect -971 -383 -925 -336
rect -971 -417 -965 -383
rect -931 -417 -925 -383
rect -971 -455 -925 -417
rect -971 -489 -965 -455
rect -931 -489 -925 -455
rect -971 -536 -925 -489
rect -813 -383 -767 -336
rect -813 -417 -807 -383
rect -773 -417 -767 -383
rect -813 -455 -767 -417
rect -813 -489 -807 -455
rect -773 -489 -767 -455
rect -813 -536 -767 -489
rect -655 -383 -609 -336
rect -655 -417 -649 -383
rect -615 -417 -609 -383
rect -655 -455 -609 -417
rect -655 -489 -649 -455
rect -615 -489 -609 -455
rect -655 -536 -609 -489
rect -497 -383 -451 -336
rect -497 -417 -491 -383
rect -457 -417 -451 -383
rect -497 -455 -451 -417
rect -497 -489 -491 -455
rect -457 -489 -451 -455
rect -497 -536 -451 -489
rect -339 -383 -293 -336
rect -339 -417 -333 -383
rect -299 -417 -293 -383
rect -339 -455 -293 -417
rect -339 -489 -333 -455
rect -299 -489 -293 -455
rect -339 -536 -293 -489
rect -181 -383 -135 -336
rect -181 -417 -175 -383
rect -141 -417 -135 -383
rect -181 -455 -135 -417
rect -181 -489 -175 -455
rect -141 -489 -135 -455
rect -181 -536 -135 -489
rect -23 -383 23 -336
rect -23 -417 -17 -383
rect 17 -417 23 -383
rect -23 -455 23 -417
rect -23 -489 -17 -455
rect 17 -489 23 -455
rect -23 -536 23 -489
rect 135 -383 181 -336
rect 135 -417 141 -383
rect 175 -417 181 -383
rect 135 -455 181 -417
rect 135 -489 141 -455
rect 175 -489 181 -455
rect 135 -536 181 -489
rect 293 -383 339 -336
rect 293 -417 299 -383
rect 333 -417 339 -383
rect 293 -455 339 -417
rect 293 -489 299 -455
rect 333 -489 339 -455
rect 293 -536 339 -489
rect 451 -383 497 -336
rect 451 -417 457 -383
rect 491 -417 497 -383
rect 451 -455 497 -417
rect 451 -489 457 -455
rect 491 -489 497 -455
rect 451 -536 497 -489
rect 609 -383 655 -336
rect 609 -417 615 -383
rect 649 -417 655 -383
rect 609 -455 655 -417
rect 609 -489 615 -455
rect 649 -489 655 -455
rect 609 -536 655 -489
rect 767 -383 813 -336
rect 767 -417 773 -383
rect 807 -417 813 -383
rect 767 -455 813 -417
rect 767 -489 773 -455
rect 807 -489 813 -455
rect 767 -536 813 -489
rect 925 -383 971 -336
rect 925 -417 931 -383
rect 965 -417 971 -383
rect 925 -455 971 -417
rect 925 -489 931 -455
rect 965 -489 971 -455
rect 925 -536 971 -489
rect 1083 -383 1129 -336
rect 1083 -417 1089 -383
rect 1123 -417 1129 -383
rect 1083 -455 1129 -417
rect 1083 -489 1089 -455
rect 1123 -489 1129 -455
rect 1083 -536 1129 -489
rect 1241 -383 1287 -336
rect 1241 -417 1247 -383
rect 1281 -417 1287 -383
rect 1241 -455 1287 -417
rect 1241 -489 1247 -455
rect 1281 -489 1287 -455
rect 1241 -536 1287 -489
rect 1399 -383 1445 -336
rect 1399 -417 1405 -383
rect 1439 -417 1445 -383
rect 1399 -455 1445 -417
rect 1399 -489 1405 -455
rect 1439 -489 1445 -455
rect 1399 -536 1445 -489
rect 1557 -383 1603 -336
rect 1557 -417 1563 -383
rect 1597 -417 1603 -383
rect 1557 -455 1603 -417
rect 1557 -489 1563 -455
rect 1597 -489 1603 -455
rect 1557 -536 1603 -489
rect 1715 -383 1761 -336
rect 1715 -417 1721 -383
rect 1755 -417 1761 -383
rect 1715 -455 1761 -417
rect 1715 -489 1721 -455
rect 1755 -489 1761 -455
rect 1715 -536 1761 -489
rect 1873 -383 1919 -336
rect 1873 -417 1879 -383
rect 1913 -417 1919 -383
rect 1873 -455 1919 -417
rect 1873 -489 1879 -455
rect 1913 -489 1919 -455
rect 1873 -536 1919 -489
rect 2031 -383 2077 -336
rect 2031 -417 2037 -383
rect 2071 -417 2077 -383
rect 2031 -455 2077 -417
rect 2031 -489 2037 -455
rect 2071 -489 2077 -455
rect 2031 -536 2077 -489
rect 2189 -383 2235 -336
rect 2189 -417 2195 -383
rect 2229 -417 2235 -383
rect 2189 -455 2235 -417
rect 2189 -489 2195 -455
rect 2229 -489 2235 -455
rect 2189 -536 2235 -489
rect 2347 -383 2393 -336
rect 2347 -417 2353 -383
rect 2387 -417 2393 -383
rect 2347 -455 2393 -417
rect 2347 -489 2353 -455
rect 2387 -489 2393 -455
rect 2347 -536 2393 -489
rect 2505 -383 2551 -336
rect 2505 -417 2511 -383
rect 2545 -417 2551 -383
rect 2505 -455 2551 -417
rect 2505 -489 2511 -455
rect 2545 -489 2551 -455
rect 2505 -536 2551 -489
rect 2663 -383 2709 -336
rect 2663 -417 2669 -383
rect 2703 -417 2709 -383
rect 2663 -455 2709 -417
rect 2663 -489 2669 -455
rect 2703 -489 2709 -455
rect 2663 -536 2709 -489
rect 2821 -383 2867 -336
rect 2821 -417 2827 -383
rect 2861 -417 2867 -383
rect 2821 -455 2867 -417
rect 2821 -489 2827 -455
rect 2861 -489 2867 -455
rect 2821 -536 2867 -489
rect 2979 -383 3025 -336
rect 2979 -417 2985 -383
rect 3019 -417 3025 -383
rect 2979 -455 3025 -417
rect 2979 -489 2985 -455
rect 3019 -489 3025 -455
rect 2979 -536 3025 -489
rect 3137 -383 3183 -336
rect 3137 -417 3143 -383
rect 3177 -417 3183 -383
rect 3137 -455 3183 -417
rect 3137 -489 3143 -455
rect 3177 -489 3183 -455
rect 3137 -536 3183 -489
rect -3127 -583 -3035 -577
rect -3127 -617 -3098 -583
rect -3064 -617 -3035 -583
rect -3127 -623 -3035 -617
rect -2969 -583 -2877 -577
rect -2969 -617 -2940 -583
rect -2906 -617 -2877 -583
rect -2969 -623 -2877 -617
rect -2811 -583 -2719 -577
rect -2811 -617 -2782 -583
rect -2748 -617 -2719 -583
rect -2811 -623 -2719 -617
rect -2653 -583 -2561 -577
rect -2653 -617 -2624 -583
rect -2590 -617 -2561 -583
rect -2653 -623 -2561 -617
rect -2495 -583 -2403 -577
rect -2495 -617 -2466 -583
rect -2432 -617 -2403 -583
rect -2495 -623 -2403 -617
rect -2337 -583 -2245 -577
rect -2337 -617 -2308 -583
rect -2274 -617 -2245 -583
rect -2337 -623 -2245 -617
rect -2179 -583 -2087 -577
rect -2179 -617 -2150 -583
rect -2116 -617 -2087 -583
rect -2179 -623 -2087 -617
rect -2021 -583 -1929 -577
rect -2021 -617 -1992 -583
rect -1958 -617 -1929 -583
rect -2021 -623 -1929 -617
rect -1863 -583 -1771 -577
rect -1863 -617 -1834 -583
rect -1800 -617 -1771 -583
rect -1863 -623 -1771 -617
rect -1705 -583 -1613 -577
rect -1705 -617 -1676 -583
rect -1642 -617 -1613 -583
rect -1705 -623 -1613 -617
rect -1547 -583 -1455 -577
rect -1547 -617 -1518 -583
rect -1484 -617 -1455 -583
rect -1547 -623 -1455 -617
rect -1389 -583 -1297 -577
rect -1389 -617 -1360 -583
rect -1326 -617 -1297 -583
rect -1389 -623 -1297 -617
rect -1231 -583 -1139 -577
rect -1231 -617 -1202 -583
rect -1168 -617 -1139 -583
rect -1231 -623 -1139 -617
rect -1073 -583 -981 -577
rect -1073 -617 -1044 -583
rect -1010 -617 -981 -583
rect -1073 -623 -981 -617
rect -915 -583 -823 -577
rect -915 -617 -886 -583
rect -852 -617 -823 -583
rect -915 -623 -823 -617
rect -757 -583 -665 -577
rect -757 -617 -728 -583
rect -694 -617 -665 -583
rect -757 -623 -665 -617
rect -599 -583 -507 -577
rect -599 -617 -570 -583
rect -536 -617 -507 -583
rect -599 -623 -507 -617
rect -441 -583 -349 -577
rect -441 -617 -412 -583
rect -378 -617 -349 -583
rect -441 -623 -349 -617
rect -283 -583 -191 -577
rect -283 -617 -254 -583
rect -220 -617 -191 -583
rect -283 -623 -191 -617
rect -125 -583 -33 -577
rect -125 -617 -96 -583
rect -62 -617 -33 -583
rect -125 -623 -33 -617
rect 33 -583 125 -577
rect 33 -617 62 -583
rect 96 -617 125 -583
rect 33 -623 125 -617
rect 191 -583 283 -577
rect 191 -617 220 -583
rect 254 -617 283 -583
rect 191 -623 283 -617
rect 349 -583 441 -577
rect 349 -617 378 -583
rect 412 -617 441 -583
rect 349 -623 441 -617
rect 507 -583 599 -577
rect 507 -617 536 -583
rect 570 -617 599 -583
rect 507 -623 599 -617
rect 665 -583 757 -577
rect 665 -617 694 -583
rect 728 -617 757 -583
rect 665 -623 757 -617
rect 823 -583 915 -577
rect 823 -617 852 -583
rect 886 -617 915 -583
rect 823 -623 915 -617
rect 981 -583 1073 -577
rect 981 -617 1010 -583
rect 1044 -617 1073 -583
rect 981 -623 1073 -617
rect 1139 -583 1231 -577
rect 1139 -617 1168 -583
rect 1202 -617 1231 -583
rect 1139 -623 1231 -617
rect 1297 -583 1389 -577
rect 1297 -617 1326 -583
rect 1360 -617 1389 -583
rect 1297 -623 1389 -617
rect 1455 -583 1547 -577
rect 1455 -617 1484 -583
rect 1518 -617 1547 -583
rect 1455 -623 1547 -617
rect 1613 -583 1705 -577
rect 1613 -617 1642 -583
rect 1676 -617 1705 -583
rect 1613 -623 1705 -617
rect 1771 -583 1863 -577
rect 1771 -617 1800 -583
rect 1834 -617 1863 -583
rect 1771 -623 1863 -617
rect 1929 -583 2021 -577
rect 1929 -617 1958 -583
rect 1992 -617 2021 -583
rect 1929 -623 2021 -617
rect 2087 -583 2179 -577
rect 2087 -617 2116 -583
rect 2150 -617 2179 -583
rect 2087 -623 2179 -617
rect 2245 -583 2337 -577
rect 2245 -617 2274 -583
rect 2308 -617 2337 -583
rect 2245 -623 2337 -617
rect 2403 -583 2495 -577
rect 2403 -617 2432 -583
rect 2466 -617 2495 -583
rect 2403 -623 2495 -617
rect 2561 -583 2653 -577
rect 2561 -617 2590 -583
rect 2624 -617 2653 -583
rect 2561 -623 2653 -617
rect 2719 -583 2811 -577
rect 2719 -617 2748 -583
rect 2782 -617 2811 -583
rect 2719 -623 2811 -617
rect 2877 -583 2969 -577
rect 2877 -617 2906 -583
rect 2940 -617 2969 -583
rect 2877 -623 2969 -617
rect 3035 -583 3127 -577
rect 3035 -617 3064 -583
rect 3098 -617 3127 -583
rect 3035 -623 3127 -617
rect -3127 -691 -3035 -685
rect -3127 -725 -3098 -691
rect -3064 -725 -3035 -691
rect -3127 -731 -3035 -725
rect -2969 -691 -2877 -685
rect -2969 -725 -2940 -691
rect -2906 -725 -2877 -691
rect -2969 -731 -2877 -725
rect -2811 -691 -2719 -685
rect -2811 -725 -2782 -691
rect -2748 -725 -2719 -691
rect -2811 -731 -2719 -725
rect -2653 -691 -2561 -685
rect -2653 -725 -2624 -691
rect -2590 -725 -2561 -691
rect -2653 -731 -2561 -725
rect -2495 -691 -2403 -685
rect -2495 -725 -2466 -691
rect -2432 -725 -2403 -691
rect -2495 -731 -2403 -725
rect -2337 -691 -2245 -685
rect -2337 -725 -2308 -691
rect -2274 -725 -2245 -691
rect -2337 -731 -2245 -725
rect -2179 -691 -2087 -685
rect -2179 -725 -2150 -691
rect -2116 -725 -2087 -691
rect -2179 -731 -2087 -725
rect -2021 -691 -1929 -685
rect -2021 -725 -1992 -691
rect -1958 -725 -1929 -691
rect -2021 -731 -1929 -725
rect -1863 -691 -1771 -685
rect -1863 -725 -1834 -691
rect -1800 -725 -1771 -691
rect -1863 -731 -1771 -725
rect -1705 -691 -1613 -685
rect -1705 -725 -1676 -691
rect -1642 -725 -1613 -691
rect -1705 -731 -1613 -725
rect -1547 -691 -1455 -685
rect -1547 -725 -1518 -691
rect -1484 -725 -1455 -691
rect -1547 -731 -1455 -725
rect -1389 -691 -1297 -685
rect -1389 -725 -1360 -691
rect -1326 -725 -1297 -691
rect -1389 -731 -1297 -725
rect -1231 -691 -1139 -685
rect -1231 -725 -1202 -691
rect -1168 -725 -1139 -691
rect -1231 -731 -1139 -725
rect -1073 -691 -981 -685
rect -1073 -725 -1044 -691
rect -1010 -725 -981 -691
rect -1073 -731 -981 -725
rect -915 -691 -823 -685
rect -915 -725 -886 -691
rect -852 -725 -823 -691
rect -915 -731 -823 -725
rect -757 -691 -665 -685
rect -757 -725 -728 -691
rect -694 -725 -665 -691
rect -757 -731 -665 -725
rect -599 -691 -507 -685
rect -599 -725 -570 -691
rect -536 -725 -507 -691
rect -599 -731 -507 -725
rect -441 -691 -349 -685
rect -441 -725 -412 -691
rect -378 -725 -349 -691
rect -441 -731 -349 -725
rect -283 -691 -191 -685
rect -283 -725 -254 -691
rect -220 -725 -191 -691
rect -283 -731 -191 -725
rect -125 -691 -33 -685
rect -125 -725 -96 -691
rect -62 -725 -33 -691
rect -125 -731 -33 -725
rect 33 -691 125 -685
rect 33 -725 62 -691
rect 96 -725 125 -691
rect 33 -731 125 -725
rect 191 -691 283 -685
rect 191 -725 220 -691
rect 254 -725 283 -691
rect 191 -731 283 -725
rect 349 -691 441 -685
rect 349 -725 378 -691
rect 412 -725 441 -691
rect 349 -731 441 -725
rect 507 -691 599 -685
rect 507 -725 536 -691
rect 570 -725 599 -691
rect 507 -731 599 -725
rect 665 -691 757 -685
rect 665 -725 694 -691
rect 728 -725 757 -691
rect 665 -731 757 -725
rect 823 -691 915 -685
rect 823 -725 852 -691
rect 886 -725 915 -691
rect 823 -731 915 -725
rect 981 -691 1073 -685
rect 981 -725 1010 -691
rect 1044 -725 1073 -691
rect 981 -731 1073 -725
rect 1139 -691 1231 -685
rect 1139 -725 1168 -691
rect 1202 -725 1231 -691
rect 1139 -731 1231 -725
rect 1297 -691 1389 -685
rect 1297 -725 1326 -691
rect 1360 -725 1389 -691
rect 1297 -731 1389 -725
rect 1455 -691 1547 -685
rect 1455 -725 1484 -691
rect 1518 -725 1547 -691
rect 1455 -731 1547 -725
rect 1613 -691 1705 -685
rect 1613 -725 1642 -691
rect 1676 -725 1705 -691
rect 1613 -731 1705 -725
rect 1771 -691 1863 -685
rect 1771 -725 1800 -691
rect 1834 -725 1863 -691
rect 1771 -731 1863 -725
rect 1929 -691 2021 -685
rect 1929 -725 1958 -691
rect 1992 -725 2021 -691
rect 1929 -731 2021 -725
rect 2087 -691 2179 -685
rect 2087 -725 2116 -691
rect 2150 -725 2179 -691
rect 2087 -731 2179 -725
rect 2245 -691 2337 -685
rect 2245 -725 2274 -691
rect 2308 -725 2337 -691
rect 2245 -731 2337 -725
rect 2403 -691 2495 -685
rect 2403 -725 2432 -691
rect 2466 -725 2495 -691
rect 2403 -731 2495 -725
rect 2561 -691 2653 -685
rect 2561 -725 2590 -691
rect 2624 -725 2653 -691
rect 2561 -731 2653 -725
rect 2719 -691 2811 -685
rect 2719 -725 2748 -691
rect 2782 -725 2811 -691
rect 2719 -731 2811 -725
rect 2877 -691 2969 -685
rect 2877 -725 2906 -691
rect 2940 -725 2969 -691
rect 2877 -731 2969 -725
rect 3035 -691 3127 -685
rect 3035 -725 3064 -691
rect 3098 -725 3127 -691
rect 3035 -731 3127 -725
rect -3183 -819 -3137 -772
rect -3183 -853 -3177 -819
rect -3143 -853 -3137 -819
rect -3183 -891 -3137 -853
rect -3183 -925 -3177 -891
rect -3143 -925 -3137 -891
rect -3183 -972 -3137 -925
rect -3025 -819 -2979 -772
rect -3025 -853 -3019 -819
rect -2985 -853 -2979 -819
rect -3025 -891 -2979 -853
rect -3025 -925 -3019 -891
rect -2985 -925 -2979 -891
rect -3025 -972 -2979 -925
rect -2867 -819 -2821 -772
rect -2867 -853 -2861 -819
rect -2827 -853 -2821 -819
rect -2867 -891 -2821 -853
rect -2867 -925 -2861 -891
rect -2827 -925 -2821 -891
rect -2867 -972 -2821 -925
rect -2709 -819 -2663 -772
rect -2709 -853 -2703 -819
rect -2669 -853 -2663 -819
rect -2709 -891 -2663 -853
rect -2709 -925 -2703 -891
rect -2669 -925 -2663 -891
rect -2709 -972 -2663 -925
rect -2551 -819 -2505 -772
rect -2551 -853 -2545 -819
rect -2511 -853 -2505 -819
rect -2551 -891 -2505 -853
rect -2551 -925 -2545 -891
rect -2511 -925 -2505 -891
rect -2551 -972 -2505 -925
rect -2393 -819 -2347 -772
rect -2393 -853 -2387 -819
rect -2353 -853 -2347 -819
rect -2393 -891 -2347 -853
rect -2393 -925 -2387 -891
rect -2353 -925 -2347 -891
rect -2393 -972 -2347 -925
rect -2235 -819 -2189 -772
rect -2235 -853 -2229 -819
rect -2195 -853 -2189 -819
rect -2235 -891 -2189 -853
rect -2235 -925 -2229 -891
rect -2195 -925 -2189 -891
rect -2235 -972 -2189 -925
rect -2077 -819 -2031 -772
rect -2077 -853 -2071 -819
rect -2037 -853 -2031 -819
rect -2077 -891 -2031 -853
rect -2077 -925 -2071 -891
rect -2037 -925 -2031 -891
rect -2077 -972 -2031 -925
rect -1919 -819 -1873 -772
rect -1919 -853 -1913 -819
rect -1879 -853 -1873 -819
rect -1919 -891 -1873 -853
rect -1919 -925 -1913 -891
rect -1879 -925 -1873 -891
rect -1919 -972 -1873 -925
rect -1761 -819 -1715 -772
rect -1761 -853 -1755 -819
rect -1721 -853 -1715 -819
rect -1761 -891 -1715 -853
rect -1761 -925 -1755 -891
rect -1721 -925 -1715 -891
rect -1761 -972 -1715 -925
rect -1603 -819 -1557 -772
rect -1603 -853 -1597 -819
rect -1563 -853 -1557 -819
rect -1603 -891 -1557 -853
rect -1603 -925 -1597 -891
rect -1563 -925 -1557 -891
rect -1603 -972 -1557 -925
rect -1445 -819 -1399 -772
rect -1445 -853 -1439 -819
rect -1405 -853 -1399 -819
rect -1445 -891 -1399 -853
rect -1445 -925 -1439 -891
rect -1405 -925 -1399 -891
rect -1445 -972 -1399 -925
rect -1287 -819 -1241 -772
rect -1287 -853 -1281 -819
rect -1247 -853 -1241 -819
rect -1287 -891 -1241 -853
rect -1287 -925 -1281 -891
rect -1247 -925 -1241 -891
rect -1287 -972 -1241 -925
rect -1129 -819 -1083 -772
rect -1129 -853 -1123 -819
rect -1089 -853 -1083 -819
rect -1129 -891 -1083 -853
rect -1129 -925 -1123 -891
rect -1089 -925 -1083 -891
rect -1129 -972 -1083 -925
rect -971 -819 -925 -772
rect -971 -853 -965 -819
rect -931 -853 -925 -819
rect -971 -891 -925 -853
rect -971 -925 -965 -891
rect -931 -925 -925 -891
rect -971 -972 -925 -925
rect -813 -819 -767 -772
rect -813 -853 -807 -819
rect -773 -853 -767 -819
rect -813 -891 -767 -853
rect -813 -925 -807 -891
rect -773 -925 -767 -891
rect -813 -972 -767 -925
rect -655 -819 -609 -772
rect -655 -853 -649 -819
rect -615 -853 -609 -819
rect -655 -891 -609 -853
rect -655 -925 -649 -891
rect -615 -925 -609 -891
rect -655 -972 -609 -925
rect -497 -819 -451 -772
rect -497 -853 -491 -819
rect -457 -853 -451 -819
rect -497 -891 -451 -853
rect -497 -925 -491 -891
rect -457 -925 -451 -891
rect -497 -972 -451 -925
rect -339 -819 -293 -772
rect -339 -853 -333 -819
rect -299 -853 -293 -819
rect -339 -891 -293 -853
rect -339 -925 -333 -891
rect -299 -925 -293 -891
rect -339 -972 -293 -925
rect -181 -819 -135 -772
rect -181 -853 -175 -819
rect -141 -853 -135 -819
rect -181 -891 -135 -853
rect -181 -925 -175 -891
rect -141 -925 -135 -891
rect -181 -972 -135 -925
rect -23 -819 23 -772
rect -23 -853 -17 -819
rect 17 -853 23 -819
rect -23 -891 23 -853
rect -23 -925 -17 -891
rect 17 -925 23 -891
rect -23 -972 23 -925
rect 135 -819 181 -772
rect 135 -853 141 -819
rect 175 -853 181 -819
rect 135 -891 181 -853
rect 135 -925 141 -891
rect 175 -925 181 -891
rect 135 -972 181 -925
rect 293 -819 339 -772
rect 293 -853 299 -819
rect 333 -853 339 -819
rect 293 -891 339 -853
rect 293 -925 299 -891
rect 333 -925 339 -891
rect 293 -972 339 -925
rect 451 -819 497 -772
rect 451 -853 457 -819
rect 491 -853 497 -819
rect 451 -891 497 -853
rect 451 -925 457 -891
rect 491 -925 497 -891
rect 451 -972 497 -925
rect 609 -819 655 -772
rect 609 -853 615 -819
rect 649 -853 655 -819
rect 609 -891 655 -853
rect 609 -925 615 -891
rect 649 -925 655 -891
rect 609 -972 655 -925
rect 767 -819 813 -772
rect 767 -853 773 -819
rect 807 -853 813 -819
rect 767 -891 813 -853
rect 767 -925 773 -891
rect 807 -925 813 -891
rect 767 -972 813 -925
rect 925 -819 971 -772
rect 925 -853 931 -819
rect 965 -853 971 -819
rect 925 -891 971 -853
rect 925 -925 931 -891
rect 965 -925 971 -891
rect 925 -972 971 -925
rect 1083 -819 1129 -772
rect 1083 -853 1089 -819
rect 1123 -853 1129 -819
rect 1083 -891 1129 -853
rect 1083 -925 1089 -891
rect 1123 -925 1129 -891
rect 1083 -972 1129 -925
rect 1241 -819 1287 -772
rect 1241 -853 1247 -819
rect 1281 -853 1287 -819
rect 1241 -891 1287 -853
rect 1241 -925 1247 -891
rect 1281 -925 1287 -891
rect 1241 -972 1287 -925
rect 1399 -819 1445 -772
rect 1399 -853 1405 -819
rect 1439 -853 1445 -819
rect 1399 -891 1445 -853
rect 1399 -925 1405 -891
rect 1439 -925 1445 -891
rect 1399 -972 1445 -925
rect 1557 -819 1603 -772
rect 1557 -853 1563 -819
rect 1597 -853 1603 -819
rect 1557 -891 1603 -853
rect 1557 -925 1563 -891
rect 1597 -925 1603 -891
rect 1557 -972 1603 -925
rect 1715 -819 1761 -772
rect 1715 -853 1721 -819
rect 1755 -853 1761 -819
rect 1715 -891 1761 -853
rect 1715 -925 1721 -891
rect 1755 -925 1761 -891
rect 1715 -972 1761 -925
rect 1873 -819 1919 -772
rect 1873 -853 1879 -819
rect 1913 -853 1919 -819
rect 1873 -891 1919 -853
rect 1873 -925 1879 -891
rect 1913 -925 1919 -891
rect 1873 -972 1919 -925
rect 2031 -819 2077 -772
rect 2031 -853 2037 -819
rect 2071 -853 2077 -819
rect 2031 -891 2077 -853
rect 2031 -925 2037 -891
rect 2071 -925 2077 -891
rect 2031 -972 2077 -925
rect 2189 -819 2235 -772
rect 2189 -853 2195 -819
rect 2229 -853 2235 -819
rect 2189 -891 2235 -853
rect 2189 -925 2195 -891
rect 2229 -925 2235 -891
rect 2189 -972 2235 -925
rect 2347 -819 2393 -772
rect 2347 -853 2353 -819
rect 2387 -853 2393 -819
rect 2347 -891 2393 -853
rect 2347 -925 2353 -891
rect 2387 -925 2393 -891
rect 2347 -972 2393 -925
rect 2505 -819 2551 -772
rect 2505 -853 2511 -819
rect 2545 -853 2551 -819
rect 2505 -891 2551 -853
rect 2505 -925 2511 -891
rect 2545 -925 2551 -891
rect 2505 -972 2551 -925
rect 2663 -819 2709 -772
rect 2663 -853 2669 -819
rect 2703 -853 2709 -819
rect 2663 -891 2709 -853
rect 2663 -925 2669 -891
rect 2703 -925 2709 -891
rect 2663 -972 2709 -925
rect 2821 -819 2867 -772
rect 2821 -853 2827 -819
rect 2861 -853 2867 -819
rect 2821 -891 2867 -853
rect 2821 -925 2827 -891
rect 2861 -925 2867 -891
rect 2821 -972 2867 -925
rect 2979 -819 3025 -772
rect 2979 -853 2985 -819
rect 3019 -853 3025 -819
rect 2979 -891 3025 -853
rect 2979 -925 2985 -891
rect 3019 -925 3025 -891
rect 2979 -972 3025 -925
rect 3137 -819 3183 -772
rect 3137 -853 3143 -819
rect 3177 -853 3183 -819
rect 3137 -891 3183 -853
rect 3137 -925 3143 -891
rect 3177 -925 3183 -891
rect 3137 -972 3183 -925
rect -3127 -1019 -3035 -1013
rect -3127 -1053 -3098 -1019
rect -3064 -1053 -3035 -1019
rect -3127 -1059 -3035 -1053
rect -2969 -1019 -2877 -1013
rect -2969 -1053 -2940 -1019
rect -2906 -1053 -2877 -1019
rect -2969 -1059 -2877 -1053
rect -2811 -1019 -2719 -1013
rect -2811 -1053 -2782 -1019
rect -2748 -1053 -2719 -1019
rect -2811 -1059 -2719 -1053
rect -2653 -1019 -2561 -1013
rect -2653 -1053 -2624 -1019
rect -2590 -1053 -2561 -1019
rect -2653 -1059 -2561 -1053
rect -2495 -1019 -2403 -1013
rect -2495 -1053 -2466 -1019
rect -2432 -1053 -2403 -1019
rect -2495 -1059 -2403 -1053
rect -2337 -1019 -2245 -1013
rect -2337 -1053 -2308 -1019
rect -2274 -1053 -2245 -1019
rect -2337 -1059 -2245 -1053
rect -2179 -1019 -2087 -1013
rect -2179 -1053 -2150 -1019
rect -2116 -1053 -2087 -1019
rect -2179 -1059 -2087 -1053
rect -2021 -1019 -1929 -1013
rect -2021 -1053 -1992 -1019
rect -1958 -1053 -1929 -1019
rect -2021 -1059 -1929 -1053
rect -1863 -1019 -1771 -1013
rect -1863 -1053 -1834 -1019
rect -1800 -1053 -1771 -1019
rect -1863 -1059 -1771 -1053
rect -1705 -1019 -1613 -1013
rect -1705 -1053 -1676 -1019
rect -1642 -1053 -1613 -1019
rect -1705 -1059 -1613 -1053
rect -1547 -1019 -1455 -1013
rect -1547 -1053 -1518 -1019
rect -1484 -1053 -1455 -1019
rect -1547 -1059 -1455 -1053
rect -1389 -1019 -1297 -1013
rect -1389 -1053 -1360 -1019
rect -1326 -1053 -1297 -1019
rect -1389 -1059 -1297 -1053
rect -1231 -1019 -1139 -1013
rect -1231 -1053 -1202 -1019
rect -1168 -1053 -1139 -1019
rect -1231 -1059 -1139 -1053
rect -1073 -1019 -981 -1013
rect -1073 -1053 -1044 -1019
rect -1010 -1053 -981 -1019
rect -1073 -1059 -981 -1053
rect -915 -1019 -823 -1013
rect -915 -1053 -886 -1019
rect -852 -1053 -823 -1019
rect -915 -1059 -823 -1053
rect -757 -1019 -665 -1013
rect -757 -1053 -728 -1019
rect -694 -1053 -665 -1019
rect -757 -1059 -665 -1053
rect -599 -1019 -507 -1013
rect -599 -1053 -570 -1019
rect -536 -1053 -507 -1019
rect -599 -1059 -507 -1053
rect -441 -1019 -349 -1013
rect -441 -1053 -412 -1019
rect -378 -1053 -349 -1019
rect -441 -1059 -349 -1053
rect -283 -1019 -191 -1013
rect -283 -1053 -254 -1019
rect -220 -1053 -191 -1019
rect -283 -1059 -191 -1053
rect -125 -1019 -33 -1013
rect -125 -1053 -96 -1019
rect -62 -1053 -33 -1019
rect -125 -1059 -33 -1053
rect 33 -1019 125 -1013
rect 33 -1053 62 -1019
rect 96 -1053 125 -1019
rect 33 -1059 125 -1053
rect 191 -1019 283 -1013
rect 191 -1053 220 -1019
rect 254 -1053 283 -1019
rect 191 -1059 283 -1053
rect 349 -1019 441 -1013
rect 349 -1053 378 -1019
rect 412 -1053 441 -1019
rect 349 -1059 441 -1053
rect 507 -1019 599 -1013
rect 507 -1053 536 -1019
rect 570 -1053 599 -1019
rect 507 -1059 599 -1053
rect 665 -1019 757 -1013
rect 665 -1053 694 -1019
rect 728 -1053 757 -1019
rect 665 -1059 757 -1053
rect 823 -1019 915 -1013
rect 823 -1053 852 -1019
rect 886 -1053 915 -1019
rect 823 -1059 915 -1053
rect 981 -1019 1073 -1013
rect 981 -1053 1010 -1019
rect 1044 -1053 1073 -1019
rect 981 -1059 1073 -1053
rect 1139 -1019 1231 -1013
rect 1139 -1053 1168 -1019
rect 1202 -1053 1231 -1019
rect 1139 -1059 1231 -1053
rect 1297 -1019 1389 -1013
rect 1297 -1053 1326 -1019
rect 1360 -1053 1389 -1019
rect 1297 -1059 1389 -1053
rect 1455 -1019 1547 -1013
rect 1455 -1053 1484 -1019
rect 1518 -1053 1547 -1019
rect 1455 -1059 1547 -1053
rect 1613 -1019 1705 -1013
rect 1613 -1053 1642 -1019
rect 1676 -1053 1705 -1019
rect 1613 -1059 1705 -1053
rect 1771 -1019 1863 -1013
rect 1771 -1053 1800 -1019
rect 1834 -1053 1863 -1019
rect 1771 -1059 1863 -1053
rect 1929 -1019 2021 -1013
rect 1929 -1053 1958 -1019
rect 1992 -1053 2021 -1019
rect 1929 -1059 2021 -1053
rect 2087 -1019 2179 -1013
rect 2087 -1053 2116 -1019
rect 2150 -1053 2179 -1019
rect 2087 -1059 2179 -1053
rect 2245 -1019 2337 -1013
rect 2245 -1053 2274 -1019
rect 2308 -1053 2337 -1019
rect 2245 -1059 2337 -1053
rect 2403 -1019 2495 -1013
rect 2403 -1053 2432 -1019
rect 2466 -1053 2495 -1019
rect 2403 -1059 2495 -1053
rect 2561 -1019 2653 -1013
rect 2561 -1053 2590 -1019
rect 2624 -1053 2653 -1019
rect 2561 -1059 2653 -1053
rect 2719 -1019 2811 -1013
rect 2719 -1053 2748 -1019
rect 2782 -1053 2811 -1019
rect 2719 -1059 2811 -1053
rect 2877 -1019 2969 -1013
rect 2877 -1053 2906 -1019
rect 2940 -1053 2969 -1019
rect 2877 -1059 2969 -1053
rect 3035 -1019 3127 -1013
rect 3035 -1053 3064 -1019
rect 3098 -1053 3127 -1019
rect 3035 -1059 3127 -1053
<< properties >>
string FIXED_BBOX -3294 -1174 3294 1174
<< end >>
