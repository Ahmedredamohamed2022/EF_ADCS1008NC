magic
tech sky130A
magscale 1 2
timestamp 1699926577
<< nwell >>
rect 4708 1220 4990 1474
rect 4708 954 5496 1220
<< metal1 >>
rect 4944 1220 4990 1632
rect 5082 1365 5508 1392
rect 5082 1313 5109 1365
rect 5161 1313 5173 1365
rect 5225 1313 5237 1365
rect 5289 1313 5301 1365
rect 5353 1313 5365 1365
rect 5417 1313 5429 1365
rect 5481 1313 5508 1365
rect 5082 1286 5508 1313
rect 2998 1164 3170 1200
rect 2998 984 3028 1164
rect 3144 984 3170 1164
rect 2998 954 3170 984
rect 3000 952 3168 954
rect 3658 866 3942 920
rect 4944 886 4992 1220
rect 5480 900 5594 960
rect 3044 558 3300 726
rect 4918 406 5528 702
rect 4806 202 5528 406
<< via1 >>
rect 5109 1313 5161 1365
rect 5173 1313 5225 1365
rect 5237 1313 5289 1365
rect 5301 1313 5353 1365
rect 5365 1313 5417 1365
rect 5429 1313 5481 1365
rect 3028 984 3144 1164
<< metal2 >>
rect 5042 1410 5518 1412
rect 3000 1408 3162 1410
rect 3684 1408 5522 1410
rect 3000 1365 5522 1408
rect 3000 1313 5109 1365
rect 5161 1313 5173 1365
rect 5225 1313 5237 1365
rect 5289 1313 5301 1365
rect 5353 1313 5365 1365
rect 5417 1313 5429 1365
rect 5481 1313 5522 1365
rect 3000 1274 5522 1313
rect 3000 1272 4910 1274
rect 3000 1270 4760 1272
rect 5042 1270 5518 1274
rect 3000 1268 4526 1270
rect 3000 1164 3162 1268
rect 3000 984 3028 1164
rect 3144 984 3162 1164
rect 3000 952 3162 984
use invm  invm_0
timestamp 1699926577
transform 1 0 2804 0 1 226
box 2164 308 2788 1248
use lsm  lsm_0
timestamp 1699926577
transform 1 0 2766 0 1 260
box -66 -58 2206 1698
<< labels >>
flabel metal1 s 5522 926 5530 946 0 FreeSans 9304 0 0 0 h0
port 1 nsew
flabel metal1 s 3062 674 3076 714 0 FreeSans 9304 0 0 0 l0
port 2 nsew
flabel metal1 s 3674 878 3682 896 0 FreeSans 3757 0 0 0 vdd1p8
port 3 nsew
flabel metal2 s 3574 1306 3582 1324 0 FreeSans 3757 0 0 0 vdd3p3
port 4 nsew
flabel metal1 s 5156 310 5198 340 0 FreeSans 3757 0 0 0 vss1p8
port 5 nsew
<< end >>
