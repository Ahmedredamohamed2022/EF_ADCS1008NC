magic
tech sky130A
magscale 1 2
timestamp 1693827120
<< metal4 >>
rect -851 438 851 600
rect -851 202 595 438
rect 831 202 851 438
rect -851 118 851 202
rect -851 -118 595 118
rect 831 -118 851 118
rect -851 -202 851 -118
rect -851 -438 595 -202
rect 831 -438 851 -202
rect -851 -600 851 -438
<< via4 >>
rect 595 202 831 438
rect 595 -118 831 118
rect 595 -438 831 -202
<< mimcap2 >>
rect -751 438 249 500
rect -751 -438 -689 438
rect 187 -438 249 438
rect -751 -500 249 -438
<< mimcap2contact >>
rect -689 -438 187 438
<< metal5 >>
rect -735 438 233 484
rect -735 -438 -689 438
rect 187 -438 233 438
rect -735 -484 233 -438
rect 553 438 873 688
rect 553 202 595 438
rect 831 202 873 438
rect 553 118 873 202
rect 553 -118 595 118
rect 831 -118 873 118
rect 553 -202 873 -118
rect 553 -438 595 -202
rect 831 -438 873 -202
rect 553 -601 873 -438
<< properties >>
string FIXED_BBOX -851 -600 349 600
<< end >>
