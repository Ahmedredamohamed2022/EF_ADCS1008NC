magic
tech sky130A
magscale 1 2
timestamp 1699289259
<< metal1 >>
rect 1700 93408 2234 93434
rect 1700 93376 1713 93408
rect 1696 93292 1713 93376
rect 2213 93376 2234 93408
rect 2213 93292 3202 93376
rect 1696 93272 3202 93292
rect 2718 90566 3124 90591
rect 2718 90322 2735 90566
rect 3107 90322 3124 90566
rect 2718 90297 3124 90322
rect 923 89763 2280 89768
rect 923 89741 2286 89763
rect 923 89625 949 89741
rect 1513 89625 2286 89741
rect 923 89566 2286 89625
rect 2086 89563 2286 89566
rect 2332 87085 2614 87109
rect 2332 86841 2351 87085
rect 2595 86841 2614 87085
rect 2332 86817 2614 86841
rect 3928 86625 4228 86671
rect 3928 85997 3960 86625
rect 4204 85997 4228 86625
rect 3928 85937 4228 85997
rect 1702 85798 2286 85843
rect 1702 85682 1737 85798
rect 2237 85682 2286 85798
rect 1702 85645 2286 85682
rect 1724 85643 2286 85645
rect 35492 85522 35982 85530
rect 2080 85498 2286 85507
rect 1718 85464 2362 85498
rect 1718 85348 1756 85464
rect 2320 85348 2362 85464
rect 34216 85484 35982 85522
rect 21980 85430 22174 85434
rect 1718 85314 2362 85348
rect 21418 85391 22174 85430
rect 2080 85297 2286 85314
rect 21418 85275 22021 85391
rect 22137 85275 22174 85391
rect 21418 85232 22174 85275
rect 21422 85231 21554 85232
rect 34216 85176 35551 85484
rect 35923 85176 35982 85484
rect 34216 85114 35982 85176
<< via1 >>
rect 1713 93292 2213 93408
rect 2735 90322 3107 90566
rect 949 89625 1513 89741
rect 2351 86841 2595 87085
rect 3960 85997 4204 86625
rect 1737 85682 2237 85798
rect 1756 85348 2320 85464
rect 22021 85275 22137 85391
rect 35551 85176 35923 85484
<< metal2 >>
rect 5340 106018 5432 106314
rect 8738 106014 8830 106310
rect 12136 106014 12228 106310
rect 15440 106012 15532 106308
rect 18750 106018 18842 106314
rect 22126 106014 22222 106316
rect 25430 106010 25526 106312
rect 28874 106010 28965 106308
rect 28794 102044 29052 102100
rect 28794 101826 28811 102044
rect 28782 101588 28811 101826
rect 29027 101588 29052 102044
rect 28782 101526 29052 101588
rect 28782 101328 29044 101526
rect 1700 93418 2234 93434
rect 1700 93408 1735 93418
rect 2191 93408 2234 93418
rect 1700 93292 1713 93408
rect 2213 93292 2234 93408
rect 1700 93282 1735 93292
rect 2191 93282 2234 93292
rect 1700 93272 2234 93282
rect 2698 93198 3034 93208
rect 2698 93142 2717 93198
rect 2773 93142 2797 93198
rect 2853 93142 2877 93198
rect 2933 93142 2957 93198
rect 3013 93142 3034 93198
rect 2322 93019 2632 93039
rect 2322 92963 2367 93019
rect 2423 92963 2447 93019
rect 2503 92963 2527 93019
rect 2583 92963 2632 93019
rect 2322 90611 2632 92963
rect 2320 90281 2632 90611
rect 914 89751 1544 89780
rect 914 89741 963 89751
rect 1499 89741 1544 89751
rect 914 89625 949 89741
rect 1513 89625 1544 89741
rect 914 89615 963 89625
rect 1499 89615 1544 89625
rect 914 89578 1544 89615
rect 2322 87085 2632 90281
rect 2698 90927 3034 93142
rect 28822 93024 29044 101328
rect 28822 92968 28862 93024
rect 28918 92968 28942 93024
rect 28998 92968 29044 93024
rect 28822 92947 29044 92968
rect 3924 92832 4224 92876
rect 3924 92536 3965 92832
rect 4181 92536 4224 92832
rect 2698 90613 3152 90927
rect 2698 90566 3158 90613
rect 2698 90322 2735 90566
rect 3107 90322 3158 90566
rect 2698 90263 3158 90322
rect 2322 86841 2351 87085
rect 2595 86841 2632 87085
rect 2322 86812 2632 86841
rect 3924 86671 4224 92536
rect 3924 86625 4228 86671
rect 3924 85997 3960 86625
rect 4204 85997 4228 86625
rect 3924 85963 4228 85997
rect 3928 85937 4228 85963
rect 1702 85808 2286 85843
rect 1702 85798 1759 85808
rect 2215 85798 2286 85808
rect 1702 85682 1737 85798
rect 2237 85682 2286 85798
rect 1702 85672 1759 85682
rect 2215 85672 2286 85682
rect 1702 85645 2286 85672
rect 1718 85474 2362 85498
rect 1718 85464 1770 85474
rect 2306 85464 2362 85474
rect 1718 85348 1756 85464
rect 2320 85348 2362 85464
rect 35492 85484 35982 85530
rect 35492 85478 35551 85484
rect 35923 85478 35982 85484
rect 1718 85338 1770 85348
rect 2306 85338 2362 85348
rect 1718 85314 2362 85338
rect 21980 85401 22174 85434
rect 21980 85265 22011 85401
rect 22147 85265 22174 85401
rect 21980 85234 22174 85265
rect 35492 85182 35549 85478
rect 35925 85182 35982 85478
rect 35492 85176 35551 85182
rect 35923 85176 35982 85182
rect 35492 85122 35982 85176
rect 34542 82969 34718 83098
rect 34542 82833 34559 82969
rect 34695 82833 34718 82969
rect 34542 82802 34718 82833
rect 20114 80021 20726 80106
rect 20114 79565 20217 80021
rect 20593 79565 20726 80021
rect 20114 79496 20726 79565
rect 20258 78572 20522 79496
rect 24506 79064 25122 79132
rect 24506 78608 24571 79064
rect 25027 78608 25122 79064
rect 33112 78778 33664 78780
rect 20286 78244 20508 78572
rect 24506 78538 25122 78608
rect 33110 78689 33674 78778
rect 24682 78252 24898 78538
rect 33110 78313 33164 78689
rect 33620 78313 33674 78689
rect 33110 78240 33674 78313
rect 33112 78222 33664 78240
rect 33248 78122 33470 78222
<< via2 >>
rect 28811 101588 29027 102044
rect 1735 93408 2191 93418
rect 1735 93292 2191 93408
rect 1735 93282 2191 93292
rect 2717 93142 2773 93198
rect 2797 93142 2853 93198
rect 2877 93142 2933 93198
rect 2957 93142 3013 93198
rect 2367 92963 2423 93019
rect 2447 92963 2503 93019
rect 2527 92963 2583 93019
rect 963 89741 1499 89751
rect 963 89625 1499 89741
rect 963 89615 1499 89625
rect 28862 92968 28918 93024
rect 28942 92968 28998 93024
rect 3965 92536 4181 92832
rect 1759 85798 2215 85808
rect 1759 85682 2215 85798
rect 1759 85672 2215 85682
rect 1770 85464 2306 85474
rect 1770 85348 2306 85464
rect 1770 85338 2306 85348
rect 22011 85391 22147 85401
rect 22011 85275 22021 85391
rect 22021 85275 22137 85391
rect 22137 85275 22147 85391
rect 22011 85265 22147 85275
rect 35549 85182 35551 85478
rect 35551 85182 35923 85478
rect 35923 85182 35925 85478
rect 34559 82833 34695 82969
rect 20217 79565 20593 80021
rect 24571 78608 25027 79064
rect 33164 78313 33620 78689
<< metal3 >>
rect 28794 102048 29052 102100
rect 28794 101584 28807 102048
rect 29031 101584 29052 102048
rect 28794 101526 29052 101584
rect 35824 100128 36132 100188
rect 35822 99990 36130 100050
rect 35826 99856 36134 99916
rect 22216 97590 22424 97630
rect 22216 97526 22247 97590
rect 22311 97526 22327 97590
rect 22391 97526 22424 97590
rect 22216 97478 22424 97526
rect 1700 93418 2234 93434
rect 1700 93382 1735 93418
rect 2191 93382 2234 93418
rect 1700 93318 1731 93382
rect 2195 93318 2234 93382
rect 1700 93282 1735 93318
rect 2191 93282 2234 93318
rect 1700 93272 2234 93282
rect 2122 93198 37208 93210
rect 2122 93142 2717 93198
rect 2773 93142 2797 93198
rect 2853 93142 2877 93198
rect 2933 93142 2957 93198
rect 3013 93196 37208 93198
rect 3013 93142 25570 93196
rect 2122 93132 25570 93142
rect 25634 93132 25650 93196
rect 25714 93132 25730 93196
rect 25794 93132 25810 93196
rect 25874 93194 37208 93196
rect 25874 93132 34972 93194
rect 2122 93130 34972 93132
rect 35036 93130 35052 93194
rect 35116 93130 35132 93194
rect 35196 93130 35212 93194
rect 35276 93130 37208 93194
rect 2122 93116 37208 93130
rect 2118 93032 37208 93040
rect 2116 93027 37208 93032
rect 2116 93024 35506 93027
rect 2116 93019 28862 93024
rect 2116 92963 2367 93019
rect 2423 92963 2447 93019
rect 2503 92963 2527 93019
rect 2583 92968 28862 93019
rect 28918 92968 28942 93024
rect 28998 92968 35506 93024
rect 2583 92963 35506 92968
rect 35570 92963 35586 93027
rect 35650 92963 35666 93027
rect 35730 92963 35746 93027
rect 35810 92963 35826 93027
rect 35890 92963 35906 93027
rect 35970 92963 37208 93027
rect 2116 92946 37208 92963
rect 2116 92942 2414 92946
rect 2116 92876 3266 92878
rect 2112 92848 37208 92876
rect 2112 92832 36159 92848
rect 2112 92536 3965 92832
rect 4181 92831 36159 92832
rect 4181 92687 22245 92831
rect 22389 92687 36159 92831
rect 4181 92544 36159 92687
rect 36543 92544 37208 92848
rect 4181 92536 37208 92544
rect 2112 92476 37208 92536
rect 2122 92354 37208 92394
rect 2122 92084 3181 92354
rect 2136 92050 3181 92084
rect 3485 92346 37208 92354
rect 3485 92050 33588 92346
rect 2136 92042 33588 92050
rect 33732 92339 37208 92346
rect 33732 92042 36757 92339
rect 2136 92035 36757 92042
rect 37141 92035 37208 92339
rect 2136 91994 37208 92035
rect 914 89751 1544 89768
rect 914 89615 963 89751
rect 1499 89615 1544 89751
rect 914 89566 1544 89615
rect 34522 86060 35334 86116
rect 1702 85812 2286 85843
rect 1702 85668 1755 85812
rect 2219 85668 2286 85812
rect 1702 85645 2286 85668
rect 34522 85676 34976 86060
rect 35280 85676 35334 86060
rect 34522 85612 35334 85676
rect 914 85500 1472 85506
rect 912 85498 2358 85500
rect 912 85478 2362 85498
rect 912 85334 1766 85478
rect 2310 85334 2362 85478
rect 35492 85482 35982 85530
rect 912 85320 2362 85334
rect 1718 85314 2362 85320
rect 21980 85401 22172 85450
rect 21980 85265 22011 85401
rect 22147 85265 22172 85401
rect 21980 83738 22172 85265
rect 35492 85178 35545 85482
rect 35929 85178 35982 85482
rect 35492 85122 35982 85178
rect 35710 85016 36124 85020
rect 33916 84824 36124 85016
rect 35710 84822 36124 84824
rect 20114 80021 20726 80106
rect 20114 79565 20217 80021
rect 20593 79904 20726 80021
rect 21982 79904 22174 83637
rect 34542 83069 34718 83098
rect 34542 82845 34555 83069
rect 34699 82845 34718 83069
rect 34542 82833 34559 82845
rect 34695 82833 34718 82845
rect 34542 82802 34718 82833
rect 20593 79712 22174 79904
rect 20593 79565 20726 79712
rect 20114 79496 20726 79565
rect 24506 79120 25122 79132
rect 1714 79116 34402 79120
rect 1714 79087 34752 79116
rect 1714 78943 1766 79087
rect 2070 79064 34752 79087
rect 2070 78943 24571 79064
rect 1714 78924 24571 78943
rect 1718 78920 24571 78924
rect 24506 78608 24571 78920
rect 25027 79045 34752 79064
rect 25027 78981 34360 79045
rect 34424 78981 34440 79045
rect 34504 78981 34520 79045
rect 34584 78981 34600 79045
rect 34664 78981 34680 79045
rect 34744 78981 34752 79045
rect 25027 78920 34752 78981
rect 25027 78608 25122 78920
rect 34322 78906 34752 78920
rect 33112 78778 33664 78780
rect 24506 78538 25122 78608
rect 33110 78689 33674 78778
rect 1716 78418 2536 78428
rect 33110 78418 33164 78689
rect 1716 78313 33164 78418
rect 33620 78313 33674 78689
rect 1716 78240 33674 78313
rect 1716 78226 33664 78240
rect 33112 78222 33664 78226
rect 34960 78016 35286 78036
rect 34960 77552 34971 78016
rect 35275 77552 35286 78016
rect 34960 77532 35286 77552
rect 35510 77233 35942 77234
rect 35510 76769 35534 77233
rect 35918 76769 35942 77233
rect 35510 76768 35942 76769
rect 36170 76411 36576 76416
rect 36170 75947 36181 76411
rect 36565 75947 36576 76411
rect 36170 75942 36576 75947
rect 36738 75608 37158 75636
rect 36738 75144 36756 75608
rect 37140 75144 37158 75608
rect 36738 75116 37158 75144
rect 2116 66716 3268 66892
rect 2120 59990 3272 60166
rect 2112 53274 3264 53450
rect 2124 46580 3276 46756
rect 2128 39810 3280 39986
rect 2116 38898 3268 39074
rect 2106 38432 3258 38608
rect 2116 32824 3268 33000
rect 2124 26118 3276 26294
rect 2120 19398 3272 19574
rect 2112 12696 3264 12872
rect 2116 5918 3268 6094
rect 2124 4378 3562 4776
rect 2118 3844 3556 4242
rect 2140 3352 3600 3740
rect 2116 2800 3598 3180
<< via3 >>
rect 28807 102044 29031 102048
rect 28807 101588 28811 102044
rect 28811 101588 29027 102044
rect 29027 101588 29031 102044
rect 28807 101584 29031 101588
rect 22247 97526 22311 97590
rect 22327 97526 22391 97590
rect 1731 93318 1735 93382
rect 1735 93318 1795 93382
rect 1811 93318 1875 93382
rect 1891 93318 1955 93382
rect 1971 93318 2035 93382
rect 2051 93318 2115 93382
rect 2131 93318 2191 93382
rect 2191 93318 2195 93382
rect 25570 93132 25634 93196
rect 25650 93132 25714 93196
rect 25730 93132 25794 93196
rect 25810 93132 25874 93196
rect 34972 93130 35036 93194
rect 35052 93130 35116 93194
rect 35132 93130 35196 93194
rect 35212 93130 35276 93194
rect 35506 92963 35570 93027
rect 35586 92963 35650 93027
rect 35666 92963 35730 93027
rect 35746 92963 35810 93027
rect 35826 92963 35890 93027
rect 35906 92963 35970 93027
rect 22245 92687 22389 92831
rect 36159 92544 36543 92848
rect 3181 92050 3485 92354
rect 33588 92042 33732 92346
rect 36757 92035 37141 92339
rect 1755 85808 2219 85812
rect 1755 85672 1759 85808
rect 1759 85672 2215 85808
rect 2215 85672 2219 85808
rect 1755 85668 2219 85672
rect 34976 85676 35280 86060
rect 1766 85474 2310 85478
rect 1766 85338 1770 85474
rect 1770 85338 2306 85474
rect 2306 85338 2310 85474
rect 1766 85334 2310 85338
rect 35545 85478 35929 85482
rect 35545 85182 35549 85478
rect 35549 85182 35925 85478
rect 35925 85182 35929 85478
rect 35545 85178 35929 85182
rect 34555 82969 34699 83069
rect 34555 82845 34559 82969
rect 34559 82845 34695 82969
rect 34695 82845 34699 82969
rect 1766 78943 2070 79087
rect 34360 78981 34424 79045
rect 34440 78981 34504 79045
rect 34520 78981 34584 79045
rect 34600 78981 34664 79045
rect 34680 78981 34744 79045
rect 34971 77552 35275 78016
rect 35534 76769 35918 77233
rect 36181 75947 36565 76411
rect 36756 75144 37140 75608
<< metal4 >>
rect 28806 102048 29032 102082
rect 28806 101584 28807 102048
rect 29031 101584 29032 102048
rect 28806 101550 29032 101584
rect 22216 97590 22424 97630
rect 22216 97526 22247 97590
rect 22311 97526 22327 97590
rect 22391 97526 22424 97590
rect 22216 97478 22424 97526
rect 1700 93382 2234 93434
rect 1700 93318 1731 93382
rect 1795 93318 1811 93382
rect 1875 93318 1891 93382
rect 1955 93318 1971 93382
rect 2035 93318 2051 93382
rect 2115 93318 2131 93382
rect 2195 93318 2234 93382
rect 1700 93272 2234 93318
rect 1704 86603 1904 93272
rect 22216 92831 22422 97478
rect 25562 93196 25882 101292
rect 25562 93132 25570 93196
rect 25634 93132 25650 93196
rect 25714 93132 25730 93196
rect 25794 93132 25810 93196
rect 25874 93132 25882 93196
rect 25562 93118 25882 93132
rect 34928 93194 35324 93208
rect 34928 93130 34972 93194
rect 35036 93130 35052 93194
rect 35116 93130 35132 93194
rect 35196 93130 35212 93194
rect 35276 93130 35324 93194
rect 22216 92687 22245 92831
rect 22389 92687 22422 92831
rect 3114 92354 3538 92394
rect 3114 92050 3181 92354
rect 3485 92050 3538 92354
rect 3114 91699 3538 92050
rect 3114 91426 3540 91699
rect 3120 91069 3540 91426
rect 22216 90497 22422 92687
rect 33539 92346 33773 92393
rect 33539 92042 33588 92346
rect 33732 92042 33773 92346
rect 33539 90477 33773 92042
rect 1688 86177 1904 86603
rect 1704 85843 1904 86177
rect 34928 86132 35324 93130
rect 35500 93027 35978 93217
rect 35500 92963 35506 93027
rect 35570 92963 35586 93027
rect 35650 92963 35666 93027
rect 35730 92963 35746 93027
rect 35810 92963 35826 93027
rect 35890 92963 35906 93027
rect 35970 92963 35978 93027
rect 34928 86060 35340 86132
rect 1702 85812 2286 85843
rect 1702 85668 1755 85812
rect 2219 85668 2286 85812
rect 1702 85645 2286 85668
rect 34928 85676 34976 86060
rect 35280 85676 35340 86060
rect 1704 85643 2284 85645
rect 1704 85641 1904 85643
rect 34928 85600 35340 85676
rect 1716 85498 1924 85504
rect 1716 85478 2362 85498
rect 1716 85334 1766 85478
rect 2310 85334 2362 85478
rect 1716 85314 2362 85334
rect 1716 79120 1924 85314
rect 34542 83069 34722 83100
rect 34542 82845 34555 83069
rect 34699 82845 34722 83069
rect 34542 82802 34722 82845
rect 1714 79087 2128 79120
rect 34542 79116 34720 82802
rect 1714 78943 1766 79087
rect 2070 78943 2128 79087
rect 1714 78924 2128 78943
rect 34322 79045 34752 79116
rect 34322 78981 34360 79045
rect 34424 78981 34440 79045
rect 34504 78981 34520 79045
rect 34584 78981 34600 79045
rect 34664 78981 34680 79045
rect 34744 78981 34752 79045
rect 34322 78906 34752 78981
rect 34928 78016 35324 85600
rect 34928 77552 34971 78016
rect 35275 77552 35324 78016
rect 34928 77466 35324 77552
rect 35500 85534 35978 92963
rect 36116 92848 36594 93209
rect 36116 92544 36159 92848
rect 36543 92544 36594 92848
rect 35500 85482 35982 85534
rect 35500 85178 35545 85482
rect 35929 85178 35982 85482
rect 35500 85122 35982 85178
rect 35500 77233 35978 85122
rect 35500 76769 35534 77233
rect 35918 76769 35978 77233
rect 35500 76695 35978 76769
rect 36116 76411 36594 92544
rect 36116 75947 36181 76411
rect 36565 75947 36594 76411
rect 36116 75897 36594 75947
rect 36718 92339 37196 93212
rect 36718 92035 36757 92339
rect 37141 92035 37196 92339
rect 36718 75608 37196 92035
rect 36718 75144 36756 75608
rect 37140 75144 37196 75608
rect 36718 75095 37196 75144
use EF_AMUX0801WISO  EF_AMUX0801WISO_0
timestamp 1699118715
transform 1 0 2428 0 -1 104312
box -306 -2006 33704 11044
use EF_DACSCA1001  EF_DACSCA1001_0
timestamp 1699118715
transform 1 0 3068 0 1 9883
box -946 -9883 66618 68998
use EF_R2RVCE  EF_R2RVCE_0
timestamp 1699118715
transform 1 0 22784 0 1 80707
box -804 -1465 11921 11144
use sample_and_hold  sample_and_hold_0
timestamp 1699118715
transform 1 0 2086 0 1 80657
box 0 -114 19469 11183
<< labels >>
flabel metal3 s 35824 100128 36132 100188 0 FreeSans 75 0 0 0 B[0]
port 1 nsew
flabel metal3 s 35822 99990 36130 100050 0 FreeSans 75 0 0 0 B[1]
port 2 nsew
flabel metal3 s 35826 99856 36134 99916 0 FreeSans 75 0 0 0 B[2]
port 3 nsew
flabel metal2 s 28874 106010 28965 106308 0 FreeSans 75 0 0 0 VIN[0]
port 4 nsew
flabel metal2 s 25430 106010 25526 106312 0 FreeSans 75 0 0 0 VIN[1]
port 5 nsew
flabel metal2 s 22126 106014 22222 106316 0 FreeSans 75 0 0 0 VIN[2]
port 6 nsew
flabel metal2 s 18750 106018 18842 106314 0 FreeSans 75 0 0 0 VIN[3]
port 7 nsew
flabel metal2 s 15440 106012 15532 106308 0 FreeSans 75 0 0 0 VIN[4]
port 8 nsew
flabel metal2 s 12136 106014 12228 106310 0 FreeSans 75 0 0 0 VIN[5]
port 9 nsew
flabel metal2 s 8738 106014 8830 106310 0 FreeSans 75 0 0 0 VIN[6]
port 10 nsew
flabel metal2 s 5340 106018 5432 106314 0 FreeSans 75 0 0 0 VIN[7]
port 11 nsew
flabel metal1 s 2086 89563 2286 89763 0 FreeSans 75 0 0 0 HOLD
port 12 nsew
flabel metal3 s 914 89566 1544 89768 0 FreeSans 4883 0 0 0 HOLD
port 12 nsew
flabel metal3 s 35710 84822 36124 85020 0 FreeSans 294 0 0 0 CMP
port 13 nsew
flabel metal3 s 2116 66716 3268 66892 0 FreeSans 6104 0 0 0 DATA[9]
port 14 nsew
flabel metal3 s 2120 59990 3272 60166 0 FreeSans 6104 0 0 0 DATA[8]
port 15 nsew
flabel metal3 s 2112 53274 3264 53450 0 FreeSans 6104 0 0 0 DATA[7]
port 16 nsew
flabel metal3 s 2124 46580 3276 46756 0 FreeSans 6104 0 0 0 DATA[6]
port 17 nsew
flabel metal3 s 2128 39810 3280 39986 0 FreeSans 6104 0 0 0 DATA[5]
port 18 nsew
flabel metal3 s 2116 32824 3268 33000 0 FreeSans 6104 0 0 0 DATA[0]
port 19 nsew
flabel metal3 s 2124 26118 3276 26294 0 FreeSans 6104 0 0 0 DATA[1]
port 20 nsew
flabel metal3 s 2120 19398 3272 19574 0 FreeSans 6104 0 0 0 DATA[2]
port 21 nsew
flabel metal3 s 2112 12696 3264 12872 0 FreeSans 6104 0 0 0 DATA[3]
port 22 nsew
flabel metal3 s 2116 5918 3268 6094 0 FreeSans 6104 0 0 0 DATA[4]
port 23 nsew
flabel metal3 s 2116 38898 3268 39074 0 FreeSans 6104 0 0 0 VH
port 24 nsew
flabel metal3 s 2106 38432 3258 38608 0 FreeSans 6104 0 0 0 VL
port 25 nsew
flabel metal3 s 1716 78226 2536 78428 0 FreeSans 6104 0 0 0 RST
port 26 nsew
flabel metal3 s 2124 4378 3562 4776 0 FreeSans 6104 0 0 0 DVDD
port 27 nsew
flabel metal3 s 2118 3844 3556 4242 0 FreeSans 6104 0 0 0 DVSS
port 28 nsew
flabel metal3 s 2116 2800 3598 3180 0 FreeSans 3906 0 0 0 VSS
port 29 nsew
flabel metal3 s 2140 3352 3600 3740 0 FreeSans 3906 0 0 0 VDD
port 30 nsew
flabel metal3 s 914 85320 1472 85506 0 FreeSans 3906 0 0 0 EN
port 31 nsew
<< end >>
