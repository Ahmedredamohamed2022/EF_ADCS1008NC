magic
tech sky130A
magscale 1 2
timestamp 1699284140
<< checkpaint >>
rect 4368 366233 76574 475071
<< metal1 >>
rect 7328 460901 7862 460927
rect 7328 460869 7341 460901
rect 7324 460785 7341 460869
rect 7841 460869 7862 460901
rect 7841 460785 8830 460869
rect 7324 460765 8830 460785
rect 8346 458059 8752 458084
rect 8346 457815 8363 458059
rect 8735 457815 8752 458059
rect 8346 457790 8752 457815
rect 6551 457256 7908 457261
rect 6551 457234 7914 457256
rect 6551 457118 6577 457234
rect 7141 457118 7914 457234
rect 6551 457059 7914 457118
rect 7714 457056 7914 457059
rect 7960 454578 8242 454602
rect 7960 454334 7979 454578
rect 8223 454334 8242 454578
rect 7960 454310 8242 454334
rect 9556 454118 9856 454164
rect 9556 453490 9588 454118
rect 9832 453490 9856 454118
rect 9556 453430 9856 453490
rect 7330 453291 7914 453336
rect 7330 453175 7365 453291
rect 7865 453175 7914 453291
rect 7330 453138 7914 453175
rect 7352 453136 7914 453138
rect 41120 453015 41610 453023
rect 7708 452991 7914 453000
rect 7346 452957 7990 452991
rect 7346 452841 7384 452957
rect 7948 452841 7990 452957
rect 39844 452977 41610 453015
rect 27608 452923 27802 452927
rect 7346 452807 7990 452841
rect 27046 452884 27802 452923
rect 7708 452790 7914 452807
rect 27046 452768 27649 452884
rect 27765 452768 27802 452884
rect 27046 452725 27802 452768
rect 27050 452724 27182 452725
rect 39844 452669 41179 452977
rect 41551 452669 41610 452977
rect 39844 452607 41610 452669
<< via1 >>
rect 7341 460785 7841 460901
rect 8363 457815 8735 458059
rect 6577 457118 7141 457234
rect 7979 454334 8223 454578
rect 9588 453490 9832 454118
rect 7365 453175 7865 453291
rect 7384 452841 7948 452957
rect 27649 452768 27765 452884
rect 41179 452669 41551 452977
<< metal2 >>
rect 10968 473511 11060 473807
rect 14366 473507 14458 473803
rect 17764 473507 17856 473803
rect 21068 473505 21160 473801
rect 24378 473511 24470 473807
rect 27754 473507 27850 473809
rect 31058 473503 31154 473805
rect 34502 473503 34593 473801
rect 34422 469537 34680 469593
rect 34422 469319 34439 469537
rect 34410 469081 34439 469319
rect 34655 469081 34680 469537
rect 34410 469019 34680 469081
rect 34410 468821 34672 469019
rect 7328 460911 7862 460927
rect 7328 460901 7363 460911
rect 7819 460901 7862 460911
rect 7328 460785 7341 460901
rect 7841 460785 7862 460901
rect 7328 460775 7363 460785
rect 7819 460775 7862 460785
rect 7328 460765 7862 460775
rect 8326 460691 8662 460701
rect 8326 460635 8345 460691
rect 8401 460635 8425 460691
rect 8481 460635 8505 460691
rect 8561 460635 8585 460691
rect 8641 460635 8662 460691
rect 7950 460512 8260 460532
rect 7950 460456 7995 460512
rect 8051 460456 8075 460512
rect 8131 460456 8155 460512
rect 8211 460456 8260 460512
rect 7950 458104 8260 460456
rect 7948 457774 8260 458104
rect 6542 457244 7172 457273
rect 6542 457234 6591 457244
rect 7127 457234 7172 457244
rect 6542 457118 6577 457234
rect 7141 457118 7172 457234
rect 6542 457108 6591 457118
rect 7127 457108 7172 457118
rect 6542 457071 7172 457108
rect 7950 454578 8260 457774
rect 8326 458420 8662 460635
rect 34450 460517 34672 468821
rect 34450 460461 34490 460517
rect 34546 460461 34570 460517
rect 34626 460461 34672 460517
rect 34450 460440 34672 460461
rect 9552 460325 9852 460369
rect 9552 460029 9593 460325
rect 9809 460029 9852 460325
rect 8326 458106 8780 458420
rect 8326 458059 8786 458106
rect 8326 457815 8363 458059
rect 8735 457815 8786 458059
rect 8326 457756 8786 457815
rect 7950 454334 7979 454578
rect 8223 454334 8260 454578
rect 7950 454305 8260 454334
rect 9552 454164 9852 460029
rect 9552 454118 9856 454164
rect 9552 453490 9588 454118
rect 9832 453490 9856 454118
rect 9552 453456 9856 453490
rect 9556 453430 9856 453456
rect 7330 453301 7914 453336
rect 7330 453291 7387 453301
rect 7843 453291 7914 453301
rect 7330 453175 7365 453291
rect 7865 453175 7914 453291
rect 7330 453165 7387 453175
rect 7843 453165 7914 453175
rect 7330 453138 7914 453165
rect 7346 452967 7990 452991
rect 7346 452957 7398 452967
rect 7934 452957 7990 452967
rect 7346 452841 7384 452957
rect 7948 452841 7990 452957
rect 41120 452977 41610 453023
rect 41120 452971 41179 452977
rect 41551 452971 41610 452977
rect 7346 452831 7398 452841
rect 7934 452831 7990 452841
rect 7346 452807 7990 452831
rect 27608 452894 27802 452927
rect 27608 452758 27639 452894
rect 27775 452758 27802 452894
rect 27608 452727 27802 452758
rect 41120 452675 41177 452971
rect 41553 452675 41610 452971
rect 41120 452669 41179 452675
rect 41551 452669 41610 452675
rect 41120 452615 41610 452669
rect 40170 450462 40346 450591
rect 40170 450326 40187 450462
rect 40323 450326 40346 450462
rect 40170 450295 40346 450326
rect 25742 447514 26354 447599
rect 25742 447058 25845 447514
rect 26221 447058 26354 447514
rect 25742 446989 26354 447058
rect 25886 446065 26150 446989
rect 30134 446557 30750 446625
rect 30134 446101 30199 446557
rect 30655 446101 30750 446557
rect 38740 446271 39292 446273
rect 25914 445737 26136 446065
rect 30134 446031 30750 446101
rect 38738 446182 39302 446271
rect 30310 445745 30526 446031
rect 38738 445806 38792 446182
rect 39248 445806 39302 446182
rect 38738 445733 39302 445806
rect 38740 445715 39292 445733
rect 38876 445615 39098 445715
<< via2 >>
rect 34439 469081 34655 469537
rect 7363 460901 7819 460911
rect 7363 460785 7819 460901
rect 7363 460775 7819 460785
rect 8345 460635 8401 460691
rect 8425 460635 8481 460691
rect 8505 460635 8561 460691
rect 8585 460635 8641 460691
rect 7995 460456 8051 460512
rect 8075 460456 8131 460512
rect 8155 460456 8211 460512
rect 6591 457234 7127 457244
rect 6591 457118 7127 457234
rect 6591 457108 7127 457118
rect 34490 460461 34546 460517
rect 34570 460461 34626 460517
rect 9593 460029 9809 460325
rect 7387 453291 7843 453301
rect 7387 453175 7843 453291
rect 7387 453165 7843 453175
rect 7398 452957 7934 452967
rect 7398 452841 7934 452957
rect 7398 452831 7934 452841
rect 27639 452884 27775 452894
rect 27639 452768 27649 452884
rect 27649 452768 27765 452884
rect 27765 452768 27775 452884
rect 27639 452758 27775 452768
rect 41177 452675 41179 452971
rect 41179 452675 41551 452971
rect 41551 452675 41553 452971
rect 40187 450326 40323 450462
rect 25845 447058 26221 447514
rect 30199 446101 30655 446557
rect 38792 445806 39248 446182
<< metal3 >>
rect 34422 469541 34680 469593
rect 34422 469077 34435 469541
rect 34659 469077 34680 469541
rect 34422 469019 34680 469077
rect 41452 467621 41760 467681
rect 41450 467483 41758 467543
rect 41454 467349 41762 467409
rect 27844 465083 28052 465123
rect 27844 465019 27875 465083
rect 27939 465019 27955 465083
rect 28019 465019 28052 465083
rect 27844 464971 28052 465019
rect 7328 460911 7862 460927
rect 7328 460875 7363 460911
rect 7819 460875 7862 460911
rect 7328 460811 7359 460875
rect 7823 460811 7862 460875
rect 7328 460775 7363 460811
rect 7819 460775 7862 460811
rect 7328 460765 7862 460775
rect 7750 460691 42836 460703
rect 7750 460635 8345 460691
rect 8401 460635 8425 460691
rect 8481 460635 8505 460691
rect 8561 460635 8585 460691
rect 8641 460689 42836 460691
rect 8641 460635 31198 460689
rect 7750 460625 31198 460635
rect 31262 460625 31278 460689
rect 31342 460625 31358 460689
rect 31422 460625 31438 460689
rect 31502 460687 42836 460689
rect 31502 460625 40600 460687
rect 7750 460623 40600 460625
rect 40664 460623 40680 460687
rect 40744 460623 40760 460687
rect 40824 460623 40840 460687
rect 40904 460623 42836 460687
rect 7750 460609 42836 460623
rect 7746 460525 42836 460533
rect 7744 460520 42836 460525
rect 7744 460517 41134 460520
rect 7744 460512 34490 460517
rect 7744 460456 7995 460512
rect 8051 460456 8075 460512
rect 8131 460456 8155 460512
rect 8211 460461 34490 460512
rect 34546 460461 34570 460517
rect 34626 460461 41134 460517
rect 8211 460456 41134 460461
rect 41198 460456 41214 460520
rect 41278 460456 41294 460520
rect 41358 460456 41374 460520
rect 41438 460456 41454 460520
rect 41518 460456 41534 460520
rect 41598 460456 42836 460520
rect 7744 460439 42836 460456
rect 7744 460435 8042 460439
rect 7744 460369 8894 460371
rect 7740 460341 42836 460369
rect 7740 460325 41787 460341
rect 7740 460029 9593 460325
rect 9809 460324 41787 460325
rect 9809 460180 27873 460324
rect 28017 460180 41787 460324
rect 9809 460037 41787 460180
rect 42171 460037 42836 460341
rect 9809 460029 42836 460037
rect 7740 459969 42836 460029
rect 7750 459847 42836 459887
rect 7750 459577 8809 459847
rect 7764 459543 8809 459577
rect 9113 459839 42836 459847
rect 9113 459543 39216 459839
rect 7764 459535 39216 459543
rect 39360 459832 42836 459839
rect 39360 459535 42385 459832
rect 7764 459528 42385 459535
rect 42769 459528 42836 459832
rect 7764 459487 42836 459528
rect 6542 457244 7172 457261
rect 6542 457108 6591 457244
rect 7127 457108 7172 457244
rect 6542 457059 7172 457108
rect 40150 453553 40962 453609
rect 7330 453305 7914 453336
rect 7330 453161 7383 453305
rect 7847 453161 7914 453305
rect 7330 453138 7914 453161
rect 40150 453169 40604 453553
rect 40908 453169 40962 453553
rect 40150 453105 40962 453169
rect 6542 452993 7100 452999
rect 6540 452991 7986 452993
rect 6540 452971 7990 452991
rect 6540 452827 7394 452971
rect 7938 452827 7990 452971
rect 41120 452975 41610 453023
rect 6540 452813 7990 452827
rect 7346 452807 7990 452813
rect 27608 452894 27800 452943
rect 27608 452758 27639 452894
rect 27775 452758 27800 452894
rect 27608 451231 27800 452758
rect 41120 452671 41173 452975
rect 41557 452671 41610 452975
rect 41120 452615 41610 452671
rect 41338 452509 41752 452513
rect 39544 452317 41752 452509
rect 41338 452315 41752 452317
rect 25742 447514 26354 447599
rect 25742 447058 25845 447514
rect 26221 447397 26354 447514
rect 27610 447397 27802 451130
rect 40170 450562 40346 450591
rect 40170 450338 40183 450562
rect 40327 450338 40346 450562
rect 40170 450326 40187 450338
rect 40323 450326 40346 450338
rect 40170 450295 40346 450326
rect 26221 447205 27802 447397
rect 26221 447058 26354 447205
rect 25742 446989 26354 447058
rect 30134 446613 30750 446625
rect 7342 446609 40030 446613
rect 7342 446580 40380 446609
rect 7342 446436 7394 446580
rect 7698 446557 40380 446580
rect 7698 446436 30199 446557
rect 7342 446417 30199 446436
rect 7346 446413 30199 446417
rect 30134 446101 30199 446413
rect 30655 446538 40380 446557
rect 30655 446474 39988 446538
rect 40052 446474 40068 446538
rect 40132 446474 40148 446538
rect 40212 446474 40228 446538
rect 40292 446474 40308 446538
rect 40372 446474 40380 446538
rect 30655 446413 40380 446474
rect 30655 446101 30750 446413
rect 39950 446399 40380 446413
rect 38740 446271 39292 446273
rect 30134 446031 30750 446101
rect 38738 446182 39302 446271
rect 7344 445911 8164 445921
rect 38738 445911 38792 446182
rect 7344 445806 38792 445911
rect 39248 445806 39302 446182
rect 7344 445733 39302 445806
rect 7344 445719 39292 445733
rect 38740 445715 39292 445719
rect 40588 445509 40914 445529
rect 40588 445045 40599 445509
rect 40903 445045 40914 445509
rect 40588 445025 40914 445045
rect 41138 444726 41570 444727
rect 41138 444262 41162 444726
rect 41546 444262 41570 444726
rect 41138 444261 41570 444262
rect 41798 443904 42204 443909
rect 41798 443440 41809 443904
rect 42193 443440 42204 443904
rect 41798 443435 42204 443440
rect 42366 443101 42786 443129
rect 42366 442637 42384 443101
rect 42768 442637 42786 443101
rect 42366 442609 42786 442637
rect 7744 434209 8896 434385
rect 7748 427483 8900 427659
rect 7740 420767 8892 420943
rect 7752 414073 8904 414249
rect 7756 407303 8908 407479
rect 7744 406391 8896 406567
rect 7734 405925 8886 406101
rect 7744 400317 8896 400493
rect 7752 393611 8904 393787
rect 7748 386891 8900 387067
rect 7740 380189 8892 380365
rect 7744 373411 8896 373587
rect 7752 371871 9190 372269
rect 7746 371337 9184 371735
rect 7768 370845 9228 371233
rect 7744 370293 9226 370673
<< via3 >>
rect 34435 469537 34659 469541
rect 34435 469081 34439 469537
rect 34439 469081 34655 469537
rect 34655 469081 34659 469537
rect 34435 469077 34659 469081
rect 27875 465019 27939 465083
rect 27955 465019 28019 465083
rect 7359 460811 7363 460875
rect 7363 460811 7423 460875
rect 7439 460811 7503 460875
rect 7519 460811 7583 460875
rect 7599 460811 7663 460875
rect 7679 460811 7743 460875
rect 7759 460811 7819 460875
rect 7819 460811 7823 460875
rect 31198 460625 31262 460689
rect 31278 460625 31342 460689
rect 31358 460625 31422 460689
rect 31438 460625 31502 460689
rect 40600 460623 40664 460687
rect 40680 460623 40744 460687
rect 40760 460623 40824 460687
rect 40840 460623 40904 460687
rect 41134 460456 41198 460520
rect 41214 460456 41278 460520
rect 41294 460456 41358 460520
rect 41374 460456 41438 460520
rect 41454 460456 41518 460520
rect 41534 460456 41598 460520
rect 27873 460180 28017 460324
rect 41787 460037 42171 460341
rect 8809 459543 9113 459847
rect 39216 459535 39360 459839
rect 42385 459528 42769 459832
rect 7383 453301 7847 453305
rect 7383 453165 7387 453301
rect 7387 453165 7843 453301
rect 7843 453165 7847 453301
rect 7383 453161 7847 453165
rect 40604 453169 40908 453553
rect 7394 452967 7938 452971
rect 7394 452831 7398 452967
rect 7398 452831 7934 452967
rect 7934 452831 7938 452967
rect 7394 452827 7938 452831
rect 41173 452971 41557 452975
rect 41173 452675 41177 452971
rect 41177 452675 41553 452971
rect 41553 452675 41557 452971
rect 41173 452671 41557 452675
rect 40183 450462 40327 450562
rect 40183 450338 40187 450462
rect 40187 450338 40323 450462
rect 40323 450338 40327 450462
rect 7394 446436 7698 446580
rect 39988 446474 40052 446538
rect 40068 446474 40132 446538
rect 40148 446474 40212 446538
rect 40228 446474 40292 446538
rect 40308 446474 40372 446538
rect 40599 445045 40903 445509
rect 41162 444262 41546 444726
rect 41809 443440 42193 443904
rect 42384 442637 42768 443101
<< metal4 >>
rect 34434 469541 34660 469575
rect 34434 469077 34435 469541
rect 34659 469077 34660 469541
rect 34434 469043 34660 469077
rect 27844 465083 28052 465123
rect 27844 465019 27875 465083
rect 27939 465019 27955 465083
rect 28019 465019 28052 465083
rect 27844 464971 28052 465019
rect 7328 460875 7862 460927
rect 7328 460811 7359 460875
rect 7423 460811 7439 460875
rect 7503 460811 7519 460875
rect 7583 460811 7599 460875
rect 7663 460811 7679 460875
rect 7743 460811 7759 460875
rect 7823 460811 7862 460875
rect 7328 460765 7862 460811
rect 7332 454096 7532 460765
rect 27844 460324 28050 464971
rect 31190 460689 31510 468785
rect 31190 460625 31198 460689
rect 31262 460625 31278 460689
rect 31342 460625 31358 460689
rect 31422 460625 31438 460689
rect 31502 460625 31510 460689
rect 31190 460611 31510 460625
rect 40556 460687 40952 460701
rect 40556 460623 40600 460687
rect 40664 460623 40680 460687
rect 40744 460623 40760 460687
rect 40824 460623 40840 460687
rect 40904 460623 40952 460687
rect 27844 460180 27873 460324
rect 28017 460180 28050 460324
rect 8742 459847 9166 459887
rect 8742 459543 8809 459847
rect 9113 459543 9166 459847
rect 8742 459192 9166 459543
rect 8742 458919 9168 459192
rect 8748 458562 9168 458919
rect 27844 457990 28050 460180
rect 39167 459839 39401 459886
rect 39167 459535 39216 459839
rect 39360 459535 39401 459839
rect 39167 457970 39401 459535
rect 7316 453670 7532 454096
rect 7332 453336 7532 453670
rect 40556 453625 40952 460623
rect 41128 460520 41606 460710
rect 41128 460456 41134 460520
rect 41198 460456 41214 460520
rect 41278 460456 41294 460520
rect 41358 460456 41374 460520
rect 41438 460456 41454 460520
rect 41518 460456 41534 460520
rect 41598 460456 41606 460520
rect 40556 453553 40968 453625
rect 7330 453305 7914 453336
rect 7330 453161 7383 453305
rect 7847 453161 7914 453305
rect 7330 453138 7914 453161
rect 40556 453169 40604 453553
rect 40908 453169 40968 453553
rect 7332 453136 7912 453138
rect 7332 453134 7532 453136
rect 40556 453093 40968 453169
rect 7344 452991 7552 452997
rect 7344 452971 7990 452991
rect 7344 452827 7394 452971
rect 7938 452827 7990 452971
rect 7344 452807 7990 452827
rect 7344 446613 7552 452807
rect 40170 450562 40350 450593
rect 40170 450338 40183 450562
rect 40327 450338 40350 450562
rect 40170 450295 40350 450338
rect 7342 446580 7756 446613
rect 40170 446609 40348 450295
rect 7342 446436 7394 446580
rect 7698 446436 7756 446580
rect 7342 446417 7756 446436
rect 39950 446538 40380 446609
rect 39950 446474 39988 446538
rect 40052 446474 40068 446538
rect 40132 446474 40148 446538
rect 40212 446474 40228 446538
rect 40292 446474 40308 446538
rect 40372 446474 40380 446538
rect 39950 446399 40380 446474
rect 40556 445509 40952 453093
rect 40556 445045 40599 445509
rect 40903 445045 40952 445509
rect 40556 444959 40952 445045
rect 41128 453027 41606 460456
rect 41744 460341 42222 460702
rect 41744 460037 41787 460341
rect 42171 460037 42222 460341
rect 41128 452975 41610 453027
rect 41128 452671 41173 452975
rect 41557 452671 41610 452975
rect 41128 452615 41610 452671
rect 41128 444726 41606 452615
rect 41128 444262 41162 444726
rect 41546 444262 41606 444726
rect 41128 444188 41606 444262
rect 41744 443904 42222 460037
rect 41744 443440 41809 443904
rect 42193 443440 42222 443904
rect 41744 443390 42222 443440
rect 42346 459832 42824 460705
rect 42346 459528 42385 459832
rect 42769 459528 42824 459832
rect 42346 443101 42824 459528
rect 42346 442637 42384 443101
rect 42768 442637 42824 443101
rect 42346 442588 42824 442637
use EF_AMUX0801WISO  EF_AMUX0801WISO_0
timestamp 1699118715
transform 1 0 8056 0 -1 471805
box -306 -2006 33704 11044
use EF_DACSCA1001  EF_DACSCA1001_0
timestamp 1699118715
transform 1 0 8696 0 1 377376
box -946 -9883 66618 68998
use EF_R2RVCE  EF_R2RVCE_0
timestamp 1699118715
transform 1 0 28412 0 1 448200
box -804 -1465 11921 11144
use sample_and_hold  sample_and_hold_0
timestamp 1699118715
transform 1 0 7714 0 1 448150
box 0 -114 19469 11183
<< labels >>
flabel metal3 s 41452 467621 41760 467681 0 FreeSans 75 0 0 0 B[0]
port 1 nsew
flabel metal3 s 41450 467483 41758 467543 0 FreeSans 75 0 0 0 B[1]
port 2 nsew
flabel metal3 s 41454 467349 41762 467409 0 FreeSans 75 0 0 0 B[2]
port 3 nsew
flabel metal2 s 34502 473503 34593 473801 0 FreeSans 75 0 0 0 VIN[0]
port 4 nsew
flabel metal2 s 31058 473503 31154 473805 0 FreeSans 75 0 0 0 VIN[1]
port 5 nsew
flabel metal2 s 27754 473507 27850 473809 0 FreeSans 75 0 0 0 VIN[2]
port 6 nsew
flabel metal2 s 24378 473511 24470 473807 0 FreeSans 75 0 0 0 VIN[3]
port 7 nsew
flabel metal2 s 21068 473505 21160 473801 0 FreeSans 75 0 0 0 VIN[4]
port 8 nsew
flabel metal2 s 17764 473507 17856 473803 0 FreeSans 75 0 0 0 VIN[5]
port 9 nsew
flabel metal2 s 14366 473507 14458 473803 0 FreeSans 75 0 0 0 VIN[6]
port 10 nsew
flabel metal2 s 10968 473511 11060 473807 0 FreeSans 75 0 0 0 VIN[7]
port 11 nsew
flabel metal1 s 7714 457056 7914 457256 0 FreeSans 75 0 0 0 HOLD
port 12 nsew
flabel metal3 s 6542 457059 7172 457261 0 FreeSans 4883 0 0 0 HOLD
port 12 nsew
flabel metal3 s 41338 452315 41752 452513 0 FreeSans 294 0 0 0 CMP
port 13 nsew
flabel metal3 s 7744 434209 8896 434385 0 FreeSans 6104 0 0 0 DATA[9]
port 14 nsew
flabel metal3 s 7748 427483 8900 427659 0 FreeSans 6104 0 0 0 DATA[8]
port 15 nsew
flabel metal3 s 7740 420767 8892 420943 0 FreeSans 6104 0 0 0 DATA[7]
port 16 nsew
flabel metal3 s 7752 414073 8904 414249 0 FreeSans 6104 0 0 0 DATA[6]
port 17 nsew
flabel metal3 s 7756 407303 8908 407479 0 FreeSans 6104 0 0 0 DATA[5]
port 18 nsew
flabel metal3 s 7744 400317 8896 400493 0 FreeSans 6104 0 0 0 DATA[0]
port 19 nsew
flabel metal3 s 7752 393611 8904 393787 0 FreeSans 6104 0 0 0 DATA[1]
port 20 nsew
flabel metal3 s 7748 386891 8900 387067 0 FreeSans 6104 0 0 0 DATA[2]
port 21 nsew
flabel metal3 s 7740 380189 8892 380365 0 FreeSans 6104 0 0 0 DATA[3]
port 22 nsew
flabel metal3 s 7744 373411 8896 373587 0 FreeSans 6104 0 0 0 DATA[4]
port 23 nsew
flabel metal3 s 7744 406391 8896 406567 0 FreeSans 6104 0 0 0 VH
port 24 nsew
flabel metal3 s 7734 405925 8886 406101 0 FreeSans 6104 0 0 0 VL
port 25 nsew
flabel metal3 s 7344 445719 8164 445921 0 FreeSans 6104 0 0 0 RST
port 26 nsew
flabel metal3 s 7752 371871 9190 372269 0 FreeSans 6104 0 0 0 DVDD
port 27 nsew
flabel metal3 s 7746 371337 9184 371735 0 FreeSans 6104 0 0 0 DVSS
port 28 nsew
flabel metal3 s 7744 370293 9226 370673 0 FreeSans 3906 0 0 0 VSS
port 29 nsew
flabel metal3 s 7768 370845 9228 371233 0 FreeSans 3906 0 0 0 VDD
port 30 nsew
flabel metal3 s 6542 452813 7100 452999 0 FreeSans 3906 0 0 0 EN
port 31 nsew
<< end >>
