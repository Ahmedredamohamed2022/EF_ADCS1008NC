magic
tech sky130A
magscale 1 2
timestamp 1694031861
<< metal1 >>
rect -2408 8024 -328 8086
rect -7490 8020 -328 8024
rect -7490 7840 -2344 8020
rect -372 7840 -328 8020
rect -7490 7836 -328 7840
rect -2408 7794 -328 7836
rect -2416 5330 -328 5350
rect -7524 5308 -328 5330
rect -7524 5128 -2301 5308
rect -393 5128 -328 5308
rect -7524 5114 -328 5128
rect -2416 5056 -328 5114
rect 2324 2602 4404 2632
rect -7554 2588 4404 2602
rect -7554 2472 2454 2588
rect 3210 2472 4404 2588
rect -7554 2446 4404 2472
rect 2324 2420 4404 2446
rect 2404 -228 4472 -198
rect -7616 -344 2583 -228
rect 4363 -344 4472 -228
rect -7616 -348 4472 -344
rect 2404 -382 4472 -348
rect 9590 -306 11676 -244
rect -2 -514 2068 -490
rect 9590 -514 9628 -306
rect -7587 -519 9628 -514
rect -7587 -635 40 -519
rect 2012 -614 9628 -519
rect 11600 -614 11676 -306
rect 2012 -635 11676 -614
rect -7587 -644 11676 -635
rect -2 -654 2068 -644
rect 9590 -652 11676 -644
rect 2398 -2998 4474 -2976
rect -7948 -3014 4474 -2998
rect -7948 -3130 2509 -3014
rect 4417 -3130 4474 -3014
rect -7948 -3146 4474 -3130
rect 2398 -3168 4474 -3146
rect -7760 -17360 -5042 -17172
rect -7730 -20082 -5032 -19866
rect -7718 -22750 -4992 -22594
rect -7650 -25544 -5004 -25424
rect -7958 -28326 -7502 -28196
<< via1 >>
rect -2344 7840 -372 8020
rect -2301 5128 -393 5308
rect 2454 2472 3210 2588
rect 2583 -344 4363 -228
rect 40 -635 2012 -519
rect 9628 -614 11600 -306
rect 2509 -3130 4417 -3014
<< metal2 >>
rect -2408 8020 -328 8086
rect -2408 7930 -2344 8020
rect -5004 7840 -2344 7930
rect -372 7930 -328 8020
rect 786 7930 886 8078
rect 3304 7930 3404 8084
rect 5644 7930 5744 8078
rect -372 7912 9372 7930
rect -372 7840 9460 7912
rect -5004 7830 9460 7840
rect -5004 5354 -4904 7830
rect -2408 7794 -328 7830
rect -5004 5254 -4688 5354
rect -2416 5316 -328 5350
rect 9360 5348 9460 7830
rect -2626 5308 -328 5316
rect -5004 2540 -4904 5254
rect -2626 5216 -2301 5308
rect -5004 2440 -4736 2540
rect -5004 -264 -4904 2440
rect -5004 -364 -4698 -264
rect -5004 -3030 -4904 -364
rect -5004 -3130 -4732 -3030
rect -5004 -6096 -4904 -3130
rect -2626 -3310 -2526 5216
rect -2416 5128 -2301 5216
rect -393 5128 -328 5308
rect -2416 5056 -328 5128
rect 956 5064 1056 5254
rect 4384 5222 5876 5322
rect 6686 5230 7102 5330
rect 9208 5248 9460 5348
rect 956 4964 4684 5064
rect -1512 3882 -1412 3954
rect 956 3882 1056 4964
rect -1512 3782 1056 3882
rect -1512 2436 -1412 3782
rect 2324 2588 4404 2626
rect 936 1118 1036 2536
rect 2324 2472 2454 2588
rect 3210 2472 4404 2588
rect 2324 2420 4404 2472
rect 936 1018 3454 1118
rect 970 998 1090 1018
rect 970 994 1070 998
rect 3354 -198 3454 1018
rect 2404 -228 4472 -198
rect -1474 -3074 -1374 -300
rect 2404 -344 2583 -228
rect 4363 -344 4472 -228
rect -6 -434 2068 -370
rect 2404 -382 4472 -344
rect -6 -519 2070 -434
rect -6 -598 40 -519
rect -4 -635 40 -598
rect 2012 -635 2070 -519
rect -4 -662 2070 -635
rect 3288 -1688 3388 -1650
rect 4584 -1688 4684 4964
rect 5776 2464 5876 5222
rect 5914 -1688 6014 -270
rect 3288 -1788 6014 -1688
rect 3288 -2976 3388 -1788
rect 4584 -1792 4684 -1788
rect 2398 -3014 4474 -2976
rect -1474 -3174 88 -3074
rect 2398 -3130 2509 -3014
rect 4417 -3130 4474 -3014
rect 7002 -3026 7102 5230
rect 9360 2550 9460 5248
rect 9174 2450 9460 2550
rect 9360 -230 9460 2450
rect 9188 -330 9460 -230
rect 9360 -3024 9460 -330
rect 9590 -306 11676 -244
rect 9590 -312 9628 -306
rect 11600 -312 11676 -306
rect 9590 -608 9626 -312
rect 11602 -608 11676 -312
rect 9590 -614 9628 -608
rect 11600 -614 11676 -608
rect 9590 -652 11676 -614
rect 6726 -3126 7102 -3026
rect 9170 -3124 9460 -3024
rect 2398 -3168 4474 -3130
rect -232 -3310 -132 -3174
rect 7002 -3310 7102 -3126
rect -2626 -3410 7102 -3310
rect -1474 -6096 -1374 -5912
rect 960 -6096 1060 -5902
rect 3368 -6096 3468 -5878
rect 5802 -6096 5902 -5882
rect 9316 -6096 9416 -3124
rect -5014 -6190 9416 -6096
rect -5014 -6192 9372 -6190
rect -4672 -6196 9372 -6192
<< via2 >>
rect 9626 -608 9628 -312
rect 9628 -608 11600 -312
rect 11600 -608 11602 -312
<< metal3 >>
rect -7254 10950 11660 11364
rect 3204 2442 3594 2588
rect 610 -350 1050 -222
rect 3246 -364 3680 -202
rect 5874 -368 6174 -194
rect 9590 -312 11676 -244
rect 9590 -608 9626 -312
rect 11602 -524 11676 -312
rect 11602 -608 11678 -524
rect 9590 -776 11678 -608
rect 5772 -3180 6056 -2994
rect 5720 -5932 6074 -5810
rect -7180 -8660 11688 -8262
rect -7114 -11428 -362 -10950
rect 2440 -11404 11686 -10994
<< metal4 >>
rect -6279 9338 -5845 12060
rect -4066 10918 -3622 12306
rect -1616 10918 -1172 12306
rect 886 10930 1330 12318
rect 3204 10956 3648 12344
rect 5562 10956 6006 12344
rect 8052 10984 8496 12372
rect 10476 10996 10920 12384
rect 10526 9606 10726 10996
rect -220 9432 -120 9452
rect 4566 9432 4666 9440
rect -6279 9096 -3196 9338
rect -2124 9332 6860 9432
rect 7686 9364 10736 9606
rect -6279 8332 -5845 9096
rect -7214 8120 -2738 8332
rect -6279 -4370 -5845 8120
rect -220 6688 -120 9332
rect 2134 6688 2234 9332
rect 4566 6688 4666 9332
rect 10526 8254 10726 9364
rect 7200 8124 11670 8254
rect -4006 6588 8260 6688
rect -220 3896 -120 6588
rect 2134 3896 2234 6588
rect 4566 3896 4666 6588
rect -4334 3796 9094 3896
rect -220 1114 -120 3796
rect 2134 1114 2234 3796
rect 4566 1114 4666 3796
rect -4394 1014 -118 1114
rect -220 -1704 -120 1014
rect 894 -282 1154 1102
rect 2106 1014 8540 1114
rect 2134 -1704 2234 1014
rect 4566 -1704 4666 1014
rect -4380 -1804 8716 -1704
rect -6632 -4700 -3380 -4370
rect -220 -4594 -120 -1804
rect 76 -3264 1994 -3212
rect 76 -3500 271 -3264
rect 507 -3500 591 -3264
rect 827 -3500 911 -3264
rect 1147 -3500 1231 -3264
rect 1467 -3500 1551 -3264
rect 1787 -3500 1994 -3264
rect 76 -3604 1994 -3500
rect 2134 -4594 2234 -1804
rect 4566 -4594 4666 -1804
rect 10526 -4394 10726 8124
rect -2144 -4694 6684 -4594
rect 7944 -4626 10726 -4394
rect -6279 -5684 -5845 -4700
rect -7200 -5882 -2722 -5684
rect 10526 -5756 10726 -4626
rect 7214 -5856 11678 -5756
rect -6279 -10040 -5845 -5882
rect -3878 -8626 -3434 -7238
rect -1584 -8638 -1140 -7250
rect 846 -8658 1290 -7270
rect 3204 -8606 3648 -7218
rect 10526 -7250 10726 -5856
rect 5592 -8638 6036 -7250
rect 8062 -8658 8506 -7270
rect 10420 -8638 10864 -7250
rect 92 -8793 2004 -8764
rect 92 -9029 285 -8793
rect 521 -9029 605 -8793
rect 841 -9029 925 -8793
rect 1161 -9029 1245 -8793
rect 1481 -9029 1565 -8793
rect 1801 -8810 2004 -8793
rect 1801 -9022 2006 -8810
rect 1801 -9029 2004 -9022
rect 92 -9188 2004 -9029
rect 10526 -9934 10726 -8638
rect -6279 -11419 -5772 -10040
rect -3984 -11362 -3477 -9983
rect -1570 -11388 -1063 -10009
rect -6267 -11428 -5772 -11419
rect -6 -11424 2080 -11330
rect 3166 -11374 3673 -9995
rect 5542 -11374 5986 -9986
rect 8078 -11362 8522 -9974
rect 10358 -11348 10865 -9969
rect 10526 -11356 10738 -11348
rect -6267 -14741 -5833 -11428
rect -6 -11660 101 -11424
rect 337 -11660 421 -11424
rect 657 -11660 741 -11424
rect 977 -11660 1061 -11424
rect 1297 -11660 1381 -11424
rect 1617 -11660 1701 -11424
rect 1937 -11660 2080 -11424
rect -6 -11732 2080 -11660
rect 74 -14472 1996 -14430
rect 74 -14708 272 -14472
rect 508 -14708 592 -14472
rect 828 -14708 912 -14472
rect 1148 -14708 1232 -14472
rect 1468 -14708 1552 -14472
rect 1788 -14708 1996 -14472
rect 10538 -14638 10738 -11356
rect 74 -14808 1996 -14708
rect 2136 -23058 2300 -22890
<< via4 >>
rect 271 -3500 507 -3264
rect 591 -3500 827 -3264
rect 911 -3500 1147 -3264
rect 1231 -3500 1467 -3264
rect 1551 -3500 1787 -3264
rect 285 -9029 521 -8793
rect 605 -9029 841 -8793
rect 925 -9029 1161 -8793
rect 1245 -9029 1481 -8793
rect 1565 -9029 1801 -8793
rect 101 -11660 337 -11424
rect 421 -11660 657 -11424
rect 741 -11660 977 -11424
rect 1061 -11660 1297 -11424
rect 1381 -11660 1617 -11424
rect 1701 -11660 1937 -11424
rect 272 -14708 508 -14472
rect 592 -14708 828 -14472
rect 912 -14708 1148 -14472
rect 1232 -14708 1468 -14472
rect 1552 -14708 1788 -14472
<< metal5 >>
rect 76 -3264 1994 -3212
rect 76 -3500 271 -3264
rect 507 -3500 591 -3264
rect 827 -3500 911 -3264
rect 1147 -3500 1231 -3264
rect 1467 -3500 1551 -3264
rect 1787 -3500 1994 -3264
rect 76 -3604 1994 -3500
rect 592 -8744 1216 -3604
rect 92 -8793 2002 -8744
rect 92 -9029 285 -8793
rect 521 -9029 605 -8793
rect 841 -9029 925 -8793
rect 1161 -9029 1245 -8793
rect 1481 -9029 1565 -8793
rect 1801 -9029 2002 -8793
rect 92 -9068 2002 -9029
rect -6 -11424 2080 -11330
rect -6 -11660 101 -11424
rect 337 -11660 421 -11424
rect 657 -11660 741 -11424
rect 977 -11660 1061 -11424
rect 1297 -11660 1381 -11424
rect 1617 -11660 1701 -11424
rect 1937 -11660 2080 -11424
rect -6 -11732 2080 -11660
rect 742 -14430 1202 -11732
rect 74 -14472 1996 -14430
rect 74 -14708 272 -14472
rect 508 -14708 592 -14472
rect 828 -14708 912 -14472
rect 1148 -14708 1232 -14472
rect 1468 -14708 1552 -14472
rect 1788 -14708 1996 -14472
rect 74 -14808 1996 -14708
use EF_LSB_CAP_WD  EF_LSB_CAP_WD_1
timestamp 1694031861
transform 1 0 12 0 1 -25196
box -7948 -8684 11688 13322
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_0
timestamp 1694031861
transform 0 1 8244 -1 0 906
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_1
timestamp 1694031861
transform 0 1 8238 -1 0 -1900
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_2
timestamp 1694031861
transform 0 1 3368 -1 0 3710
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_3
timestamp 1694031861
transform 0 1 10642 -1 0 -7482
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_4
timestamp 1694031861
transform 0 1 10638 -1 0 912
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_5
timestamp 1694031861
transform 0 1 3442 -1 0 902
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_6
timestamp 1694031861
transform 0 1 -6170 -1 0 3698
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_7
timestamp 1694031861
transform 0 1 1034 -1 0 3698
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_8
timestamp 1694031861
transform 0 1 10640 -1 0 3726
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_9
timestamp 1694031861
transform 0 1 10638 -1 0 6532
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_10
timestamp 1694031861
transform 0 1 10640 -1 0 9334
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_11
timestamp 1694031861
transform 0 1 10640 -1 0 -1880
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_12
timestamp 1694031861
transform 0 1 -6154 -1 0 -1886
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_13
timestamp 1694031861
transform 0 1 1030 -1 0 898
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_14
timestamp 1694031861
transform 0 1 -6168 -1 0 904
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_15
timestamp 1694031861
transform 0 1 10642 -1 0 -4684
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_16
timestamp 1694031861
transform 0 1 5840 -1 0 -7496
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_17
timestamp 1694031861
transform 0 1 5842 -1 0 904
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_18
timestamp 1694031861
transform 0 1 5842 -1 0 3706
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_19
timestamp 1694031861
transform 0 1 5838 -1 0 12116
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_20
timestamp 1694031861
transform 0 1 5842 -1 0 6508
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_21
timestamp 1694031861
transform 0 1 3436 -1 0 6500
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_22
timestamp 1694031861
transform 0 1 1034 -1 0 6500
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_23
timestamp 1694031861
transform 0 1 -6164 -1 0 6506
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_24
timestamp 1694031861
transform 0 1 -1364 -1 0 6506
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_25
timestamp 1694031861
transform 0 1 -1366 -1 0 3700
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_26
timestamp 1694031861
transform 0 1 -1368 -1 0 902
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_27
timestamp 1694031861
transform 0 1 8238 -1 0 9310
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_28
timestamp 1694031861
transform 0 1 -1362 -1 0 -1892
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_29
timestamp 1694031861
transform 0 1 1032 -1 0 -1904
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_30
timestamp 1694031861
transform 0 1 3440 -1 0 -1894
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_31
timestamp 1694031861
transform 0 1 5838 -1 0 -1898
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_32
timestamp 1694031861
transform 0 1 5844 -1 0 9312
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_33
timestamp 1694031861
transform 0 1 3440 -1 0 9302
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_34
timestamp 1694031861
transform 0 1 1036 -1 0 9302
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_35
timestamp 1694031861
transform 0 1 -6168 -1 0 12124
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_36
timestamp 1694031861
transform 0 1 -1366 -1 0 9306
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_37
timestamp 1694031861
transform 0 1 -6162 -1 0 9312
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_38
timestamp 1694031861
transform 0 1 10650 -1 0 -10208
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_39
timestamp 1694031861
transform 0 1 1034 -1 0 -7498
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_40
timestamp 1694031861
transform 0 1 3444 -1 0 -7492
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_41
timestamp 1694031861
transform 0 1 8246 -1 0 -7490
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_42
timestamp 1694031861
transform 0 1 -3764 -1 0 12118
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_43
timestamp 1694031861
transform 0 1 -3764 -1 0 9312
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_44
timestamp 1694031861
transform 0 1 -3764 -1 0 6504
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_45
timestamp 1694031861
transform 0 1 -3766 -1 0 3702
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_46
timestamp 1694031861
transform 0 1 10638 -1 0 12136
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_47
timestamp 1694031861
transform 0 1 8244 -1 0 3708
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_48
timestamp 1694031861
transform 0 1 -3764 -1 0 906
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_49
timestamp 1694031861
transform 0 1 8242 -1 0 6512
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_50
timestamp 1694031861
transform 0 1 -3760 -1 0 -1894
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_51
timestamp 1694031861
transform 0 1 -1358 -1 0 -7492
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_52
timestamp 1694031861
transform 0 1 -3756 -1 0 -7480
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_53
timestamp 1694031861
transform 0 1 8240 -1 0 12108
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_54
timestamp 1694031861
transform 0 1 3438 -1 0 12106
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_55
timestamp 1694031861
transform 0 1 1036 -1 0 12106
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_56
timestamp 1694031861
transform 0 1 8248 -1 0 -4690
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_57
timestamp 1694031861
transform 0 1 -1364 -1 0 12106
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_58
timestamp 1694031861
transform 0 1 5838 -1 0 -4696
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_59
timestamp 1694031861
transform 0 1 3442 -1 0 -4694
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_60
timestamp 1694031861
transform 0 1 1034 -1 0 -4702
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_61
timestamp 1694031861
transform 0 1 -1360 -1 0 -4690
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_62
timestamp 1694031861
transform 0 1 -3758 -1 0 -4684
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_63
timestamp 1694031861
transform 0 1 -6154 -1 0 -4680
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_64
timestamp 1694031861
transform 0 1 -6154 -1 0 -7474
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_65
timestamp 1694031861
transform 0 1 -6150 -1 0 -10260
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_66
timestamp 1694031861
transform 0 1 -3746 -1 0 -10262
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_67
timestamp 1694031861
transform 0 1 -1340 -1 0 -10252
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_68
timestamp 1694031861
transform 0 1 1052 -1 0 -10242
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_69
timestamp 1694031861
transform 0 1 3450 -1 0 -10234
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_70
timestamp 1694031861
transform 0 1 5846 -1 0 -10228
box -1186 -1040 1186 1040
use sky130_fd_pr__cap_mim_m3_1_6ZNTNB  sky130_fd_pr__cap_mim_m3_1_6ZNTNB_71
timestamp 1694031861
transform 0 1 8244 -1 0 -10222
box -1186 -1040 1186 1040
use via23  via23_0
timestamp 1694031861
transform 1 0 6875 0 1 2432
box -2079 0 1 100
use via23  via23_1
timestamp 1694031861
transform 1 0 2073 0 1 2412
box -2079 0 1 100
use via23  via23_2
timestamp 1694031861
transform 1 0 4483 0 1 -380
box -2079 0 1 100
use via23  via23_3
timestamp 1694031861
transform 1 0 2073 0 1 -382
box -2079 0 1 100
use via23  via23_4
timestamp 1694031861
transform 1 0 4481 0 1 -3172
box -2079 0 1 100
use via23  via23_5
timestamp 1694031861
transform 1 0 6879 0 1 -372
box -2079 0 1 100
use via23  via23_6
timestamp 1694031861
transform 1 0 -329 0 1 2416
box -2079 0 1 100
use via23  via23_7
timestamp 1694031861
transform 1 0 2075 0 1 5216
box -2079 0 1 100
use via23  via23_8
timestamp 1694031861
transform 1 0 2075 0 1 -3184
box -2079 0 1 100
use via23  via23_9
timestamp 1694031861
transform 1 0 -321 0 1 5226
box -2079 0 1 100
use via23  via23_10
timestamp 1694031861
transform 1 0 -329 0 1 -374
box -2079 0 1 100
use via23  via23_11
timestamp 1694031861
transform 1 0 -323 0 1 -3170
box -2079 0 1 100
use via23  via23_12
timestamp 1694031861
transform 1 0 6877 0 1 -3178
box -2079 0 1 100
use via23  via23_13
timestamp 1694031861
transform 1 0 6875 0 1 5242
box -2079 0 1 100
use via23  via23_14
timestamp 1694031861
transform 1 0 4477 0 1 5226
box -2079 0 1 100
use via23  via23_15
timestamp 1694031861
transform 1 0 4407 0 1 2424
box -2079 0 1 100
use via23  via23_16
timestamp 1694031861
transform 1 0 -325 0 1 8034
box -2079 0 1 100
use via23  via23_17
timestamp 1694031861
transform 1 0 2073 0 1 8032
box -2079 0 1 100
use via23  via23_18
timestamp 1694031861
transform 1 0 4471 0 1 8020
box -2079 0 1 100
use via23  via23_19
timestamp 1694031861
transform 1 0 9275 0 1 -3154
box -2079 0 1 100
use via23  via23_20
timestamp 1694031861
transform 1 0 6875 0 1 8032
box -2079 0 1 100
use via23  via23_21
timestamp 1694031861
transform 1 0 9275 0 1 5238
box -2079 0 1 100
use via23  via23_22
timestamp 1694031861
transform 1 0 9275 0 1 2442
box -2079 0 1 100
use via23  via23_23
timestamp 1694031861
transform 1 0 9277 0 1 -356
box -2079 0 1 100
use via23  via23_24
timestamp 1694031861
transform 1 0 -2727 0 1 -3158
box -2079 0 1 100
use via23  via23_25
timestamp 1694031861
transform 1 0 6885 0 1 -5958
box -2079 0 1 100
use via23  via23_26
timestamp 1694031861
transform 1 0 4475 0 1 -5942
box -2079 0 1 100
use via23  via23_27
timestamp 1694031861
transform 1 0 2069 0 1 -5966
box -2079 0 1 100
use via23  via23_28
timestamp 1694031861
transform 1 0 -325 0 1 -5960
box -2079 0 1 100
use via23  via23_29
timestamp 1694031861
transform 1 0 -2727 0 1 -366
box -2079 0 1 100
use via23  via23_30
timestamp 1694031861
transform 1 0 -2723 0 1 2432
box -2079 0 1 100
use via23  via23_31
timestamp 1694031861
transform 1 0 -2729 0 1 5244
box -2079 0 1 100
<< labels >>
flabel metal1 s -7490 2502 -7398 2576 0 FreeSans 1024 0 0 0 D5
port 1 nsew
flabel metal1 s -7510 -316 -7418 -242 0 FreeSans 1024 0 0 0 D6
port 2 nsew
flabel metal1 s -7730 -3106 -7638 -3032 0 FreeSans 1024 0 0 0 D7
port 3 nsew
flabel metal1 s -7482 5166 -7376 5260 0 FreeSans 1024 0 0 0 D8
port 4 nsew
flabel metal1 s -7442 7910 -7342 7998 0 FreeSans 1024 0 0 0 D9
port 5 nsew
flabel metal1 s -7496 -616 -7390 -528 0 FreeSans 1024 0 0 0 VSS
port 6 nsew
flabel metal4 s 2152 2160 2216 2320 0 FreeSans 1024 0 0 0 VP2
port 7 nsew
flabel metal4 s 2168 -23008 2232 -22944 0 FreeSans 411 0 0 0 VP1
port 8 nsew
flabel metal1 s -7668 -22694 -7542 -22604 0 FreeSans 655 0 0 0 D0
port 9 nsew
flabel metal1 s -7598 -25530 -7506 -25432 0 FreeSans 655 0 0 0 D1
port 10 nsew
flabel metal1 s -7736 -17300 -7616 -17200 0 FreeSans 655 0 0 0 D4
port 11 nsew
flabel metal1 s -7666 -20064 -7572 -19878 0 FreeSans 655 0 0 0 D3
port 12 nsew
flabel metal1 s -7678 -28290 -7610 -28248 0 FreeSans 655 0 0 0 D2
port 13 nsew
<< end >>
