magic
tech sky130A
magscale 1 2
timestamp 1699926577
<< metal1 >>
rect 12914 11016 13290 11028
rect 12914 10964 12916 11016
rect 12968 10964 12980 11016
rect 13032 10964 13044 11016
rect 13096 10964 13108 11016
rect 13160 10964 13172 11016
rect 13224 10964 13236 11016
rect 13288 10964 13290 11016
rect 12914 10952 13290 10964
rect 2746 2156 2828 2178
rect 2746 2104 2761 2156
rect 2813 2104 2828 2156
rect 2746 2092 2828 2104
rect 2746 2040 2761 2092
rect 2813 2040 2828 2092
rect 2746 2028 2828 2040
rect 2746 1976 2761 2028
rect 2813 1976 2828 2028
rect 2746 1964 2828 1976
rect 2746 1912 2761 1964
rect 2813 1912 2828 1964
rect 2746 1900 2828 1912
rect 2746 1848 2761 1900
rect 2813 1848 2828 1900
rect 2746 1826 2828 1848
rect 6112 2158 6194 2180
rect 6112 2106 6127 2158
rect 6179 2106 6194 2158
rect 6112 2094 6194 2106
rect 6112 2042 6127 2094
rect 6179 2042 6194 2094
rect 6112 2030 6194 2042
rect 6112 1978 6127 2030
rect 6179 1978 6194 2030
rect 6112 1966 6194 1978
rect 6112 1914 6127 1966
rect 6179 1914 6194 1966
rect 6112 1902 6194 1914
rect 6112 1850 6127 1902
rect 6179 1850 6194 1902
rect 6112 1828 6194 1850
rect 9462 2158 9544 2180
rect 9462 2106 9477 2158
rect 9529 2106 9544 2158
rect 9462 2094 9544 2106
rect 9462 2042 9477 2094
rect 9529 2042 9544 2094
rect 9462 2030 9544 2042
rect 9462 1978 9477 2030
rect 9529 1978 9544 2030
rect 9462 1966 9544 1978
rect 9462 1914 9477 1966
rect 9529 1914 9544 1966
rect 9462 1902 9544 1914
rect 9462 1850 9477 1902
rect 9529 1850 9544 1902
rect 9462 1828 9544 1850
rect 12834 2156 12916 2178
rect 12834 2104 12849 2156
rect 12901 2104 12916 2156
rect 12834 2092 12916 2104
rect 12834 2040 12849 2092
rect 12901 2040 12916 2092
rect 12834 2028 12916 2040
rect 12834 1976 12849 2028
rect 12901 1976 12916 2028
rect 12834 1964 12916 1976
rect 12834 1912 12849 1964
rect 12901 1912 12916 1964
rect 12834 1900 12916 1912
rect 12834 1848 12849 1900
rect 12901 1848 12916 1900
rect 12834 1826 12916 1848
rect 16130 2152 16212 2174
rect 16130 2100 16145 2152
rect 16197 2100 16212 2152
rect 16130 2088 16212 2100
rect 16130 2036 16145 2088
rect 16197 2036 16212 2088
rect 16130 2024 16212 2036
rect 16130 1972 16145 2024
rect 16197 1972 16212 2024
rect 16130 1960 16212 1972
rect 16130 1908 16145 1960
rect 16197 1908 16212 1960
rect 16130 1896 16212 1908
rect 16130 1844 16145 1896
rect 16197 1844 16212 1896
rect 16130 1822 16212 1844
rect 19506 2160 19588 2182
rect 19506 2108 19521 2160
rect 19573 2108 19588 2160
rect 19506 2096 19588 2108
rect 19506 2044 19521 2096
rect 19573 2044 19588 2096
rect 19506 2032 19588 2044
rect 19506 1980 19521 2032
rect 19573 1980 19588 2032
rect 19506 1968 19588 1980
rect 19506 1916 19521 1968
rect 19573 1916 19588 1968
rect 19506 1904 19588 1916
rect 19506 1852 19521 1904
rect 19573 1852 19588 1904
rect 19506 1830 19588 1852
rect 22852 2132 22868 2184
rect 22920 2132 22936 2184
rect 22852 2120 22936 2132
rect 22852 2068 22868 2120
rect 22920 2068 22936 2120
rect 22852 2056 22936 2068
rect 22852 2004 22868 2056
rect 22920 2004 22936 2056
rect 22852 1992 22936 2004
rect 22852 1940 22868 1992
rect 22920 1940 22936 1992
rect 22852 1928 22936 1940
rect 22852 1876 22868 1928
rect 22920 1876 22936 1928
rect 22852 1864 22936 1876
rect 22852 1812 22868 1864
rect 22920 1812 22936 1864
rect 26226 2165 26306 2192
rect 26226 2113 26240 2165
rect 26292 2113 26306 2165
rect 26226 2101 26306 2113
rect 26226 2049 26240 2101
rect 26292 2049 26306 2101
rect 26226 2037 26306 2049
rect 26226 1985 26240 2037
rect 26292 1985 26306 2037
rect 26226 1973 26306 1985
rect 26226 1921 26240 1973
rect 26292 1921 26306 1973
rect 26226 1909 26306 1921
rect 26226 1857 26240 1909
rect 26292 1857 26306 1909
rect 26226 1830 26306 1857
rect 342 494 602 522
rect 342 378 384 494
rect 564 378 602 494
rect 342 348 602 378
rect 3712 498 3974 524
rect 3712 382 3754 498
rect 3934 382 3974 498
rect 3712 348 3974 382
rect 7060 500 7324 530
rect 7060 384 7106 500
rect 7286 384 7324 500
rect 7060 348 7324 384
rect 10430 495 10696 518
rect 10430 379 10476 495
rect 10656 379 10696 495
rect 10430 356 10696 379
rect 13736 496 13986 524
rect 13736 380 13771 496
rect 13951 380 13986 496
rect 13736 350 13986 380
rect 17096 504 17364 526
rect 17096 388 17142 504
rect 17322 388 17364 504
rect 17096 356 17364 388
rect 20452 496 20718 524
rect 20452 380 20495 496
rect 20675 380 20718 496
rect 20452 346 20718 380
rect 23824 509 24082 524
rect 23824 393 23861 509
rect 24041 393 24082 509
rect 23824 362 24082 393
rect 25858 231 26306 276
rect 25858 51 25895 231
rect 26267 51 26306 231
rect 25858 8 26306 51
<< via1 >>
rect 12916 10964 12968 11016
rect 12980 10964 13032 11016
rect 13044 10964 13096 11016
rect 13108 10964 13160 11016
rect 13172 10964 13224 11016
rect 13236 10964 13288 11016
rect 2761 2104 2813 2156
rect 2761 2040 2813 2092
rect 2761 1976 2813 2028
rect 2761 1912 2813 1964
rect 2761 1848 2813 1900
rect 6127 2106 6179 2158
rect 6127 2042 6179 2094
rect 6127 1978 6179 2030
rect 6127 1914 6179 1966
rect 6127 1850 6179 1902
rect 9477 2106 9529 2158
rect 9477 2042 9529 2094
rect 9477 1978 9529 2030
rect 9477 1914 9529 1966
rect 9477 1850 9529 1902
rect 12849 2104 12901 2156
rect 12849 2040 12901 2092
rect 12849 1976 12901 2028
rect 12849 1912 12901 1964
rect 12849 1848 12901 1900
rect 16145 2100 16197 2152
rect 16145 2036 16197 2088
rect 16145 1972 16197 2024
rect 16145 1908 16197 1960
rect 16145 1844 16197 1896
rect 19521 2108 19573 2160
rect 19521 2044 19573 2096
rect 19521 1980 19573 2032
rect 19521 1916 19573 1968
rect 19521 1852 19573 1904
rect 22868 2132 22920 2184
rect 22868 2068 22920 2120
rect 22868 2004 22920 2056
rect 22868 1940 22920 1992
rect 22868 1876 22920 1928
rect 22868 1812 22920 1864
rect 26240 2113 26292 2165
rect 26240 2049 26292 2101
rect 26240 1985 26292 2037
rect 26240 1921 26292 1973
rect 26240 1857 26292 1909
rect 384 378 564 494
rect 3754 382 3934 498
rect 7106 384 7286 500
rect 10476 379 10656 495
rect 13771 380 13951 496
rect 17142 388 17322 504
rect 20495 380 20675 496
rect 23861 393 24041 509
rect 25895 51 26267 231
<< metal2 >>
rect 12900 11016 13304 11042
rect 12900 10964 12916 11016
rect 12968 10964 12980 11016
rect 13032 10964 13044 11016
rect 13096 10964 13108 11016
rect 13160 10964 13172 11016
rect 13224 10964 13236 11016
rect 13288 10964 13304 11016
rect 12900 10934 13304 10964
rect 12902 10930 13304 10934
rect 2732 2156 2836 2198
rect 2732 2104 2761 2156
rect 2813 2104 2836 2156
rect 2732 2092 2836 2104
rect 2732 2040 2761 2092
rect 2813 2040 2836 2092
rect 2732 2028 2836 2040
rect 2732 1976 2761 2028
rect 2813 2000 2836 2028
rect 6104 2158 6208 2212
rect 6104 2106 6127 2158
rect 6179 2106 6208 2158
rect 6104 2094 6208 2106
rect 6104 2042 6127 2094
rect 6179 2042 6208 2094
rect 6104 2030 6208 2042
rect 2813 1998 2920 2000
rect 2813 1976 3004 1998
rect 2732 1964 3004 1976
rect 2732 1912 2761 1964
rect 2813 1912 3004 1964
rect 2732 1906 3004 1912
rect 2732 1900 2836 1906
rect 2732 1848 2761 1900
rect 2813 1848 2836 1900
rect 2732 1800 2836 1848
rect 342 494 602 522
rect 342 378 384 494
rect 564 378 602 494
rect 56 172 228 376
rect 342 348 602 378
rect -300 154 228 172
rect -300 18 -257 154
rect -41 18 228 154
rect -300 0 228 18
rect 400 268 502 348
rect 400 -1504 494 268
rect 298 -1525 604 -1504
rect 298 -1581 336 -1525
rect 392 -1581 416 -1525
rect 472 -1581 496 -1525
rect 552 -1581 604 -1525
rect 298 -1600 604 -1581
rect 400 -1603 494 -1600
rect 2912 -1708 3004 1906
rect 6104 1978 6127 2030
rect 6179 1998 6208 2030
rect 9454 2158 9558 2200
rect 9454 2106 9477 2158
rect 9529 2106 9558 2158
rect 9454 2094 9558 2106
rect 9454 2042 9477 2094
rect 9529 2042 9558 2094
rect 9454 2030 9558 2042
rect 6179 1994 6284 1998
rect 6179 1978 6401 1994
rect 6104 1966 6401 1978
rect 6104 1914 6127 1966
rect 6179 1914 6401 1966
rect 6104 1904 6401 1914
rect 6104 1902 6208 1904
rect 6104 1850 6127 1902
rect 6179 1850 6208 1902
rect 6104 1814 6208 1850
rect 3712 498 3974 524
rect 3712 382 3754 498
rect 3934 382 3974 498
rect 3712 348 3974 382
rect 3800 288 3902 348
rect 3809 -1300 3891 288
rect 3696 -1323 4002 -1300
rect 3696 -1379 3736 -1323
rect 3792 -1379 3816 -1323
rect 3872 -1379 3896 -1323
rect 3952 -1379 4002 -1323
rect 3696 -1396 4002 -1379
rect 3809 -1397 3891 -1396
rect 2908 -2000 3004 -1708
rect 6311 -1704 6401 1904
rect 9454 1978 9477 2030
rect 9529 1998 9558 2030
rect 12828 2156 12932 2200
rect 12828 2104 12849 2156
rect 12901 2104 12932 2156
rect 12828 2092 12932 2104
rect 12828 2040 12849 2092
rect 12901 2040 12932 2092
rect 12828 2028 12932 2040
rect 9529 1994 9632 1998
rect 9529 1978 9800 1994
rect 9454 1966 9800 1978
rect 9454 1914 9477 1966
rect 9529 1914 9800 1966
rect 9454 1906 9800 1914
rect 9454 1904 9632 1906
rect 9454 1902 9558 1904
rect 9454 1850 9477 1902
rect 9529 1850 9558 1902
rect 9454 1802 9558 1850
rect 7060 500 7324 530
rect 7060 384 7106 500
rect 7286 384 7324 500
rect 7060 348 7324 384
rect 7138 280 7240 348
rect 7138 -1100 7226 280
rect 7008 -1123 7314 -1100
rect 7008 -1179 7056 -1123
rect 7112 -1179 7136 -1123
rect 7192 -1179 7216 -1123
rect 7272 -1179 7314 -1123
rect 7008 -1196 7314 -1179
rect 7138 -1198 7226 -1196
rect 9712 -1698 9800 1906
rect 12828 1976 12849 2028
rect 12901 2002 12932 2028
rect 16120 2152 16224 2206
rect 16120 2100 16145 2152
rect 16197 2100 16224 2152
rect 16120 2088 16224 2100
rect 16120 2036 16145 2088
rect 16197 2036 16224 2088
rect 16120 2024 16224 2036
rect 12901 1976 13097 2002
rect 12828 1964 13097 1976
rect 12828 1912 12849 1964
rect 12901 1912 13097 1964
rect 12828 1908 13097 1912
rect 12828 1900 12932 1908
rect 12828 1848 12849 1900
rect 12901 1848 12932 1900
rect 12828 1802 12932 1848
rect 10430 495 10696 518
rect 10430 379 10476 495
rect 10656 379 10696 495
rect 10430 356 10696 379
rect 10520 294 10622 356
rect 10532 -902 10608 294
rect 10406 -919 10712 -902
rect 10406 -975 10450 -919
rect 10506 -975 10530 -919
rect 10586 -975 10610 -919
rect 10666 -975 10712 -919
rect 10406 -998 10712 -975
rect 13019 -1698 13097 1908
rect 16120 1972 16145 2024
rect 16197 1998 16224 2024
rect 19494 2160 19598 2206
rect 19494 2108 19521 2160
rect 19573 2108 19598 2160
rect 19494 2096 19598 2108
rect 19494 2044 19521 2096
rect 19573 2044 19598 2096
rect 19494 2032 19598 2044
rect 16197 1980 16226 1998
rect 19494 1980 19521 2032
rect 19573 2004 19598 2032
rect 22840 2184 22946 2200
rect 22840 2132 22868 2184
rect 22920 2132 22946 2184
rect 22840 2120 22946 2132
rect 22840 2068 22868 2120
rect 22920 2068 22946 2120
rect 22840 2056 22946 2068
rect 22840 2004 22868 2056
rect 22920 2004 22946 2056
rect 19573 1980 19795 2004
rect 16197 1972 16400 1980
rect 16120 1960 16400 1972
rect 16120 1908 16145 1960
rect 16197 1908 16400 1960
rect 16120 1904 16400 1908
rect 16120 1896 16224 1904
rect 16120 1844 16145 1896
rect 16197 1844 16224 1896
rect 16120 1808 16224 1844
rect 13736 496 13986 524
rect 13736 380 13771 496
rect 13951 380 13986 496
rect 13736 350 13986 380
rect 13816 302 13918 350
rect 13830 -698 13898 302
rect 13706 -721 14012 -698
rect 13706 -777 13740 -721
rect 13796 -777 13820 -721
rect 13876 -777 13900 -721
rect 13956 -777 14012 -721
rect 13706 -794 14012 -777
rect 13830 -802 13898 -794
rect 2908 -2006 2998 -2000
rect 6311 -2001 6402 -1704
rect 9712 -1996 9802 -1698
rect 13012 -1996 13102 -1698
rect 16324 -1704 16400 1904
rect 19494 1968 19795 1980
rect 19494 1916 19521 1968
rect 19573 1916 19795 1968
rect 19494 1906 19795 1916
rect 19494 1904 19598 1906
rect 19494 1852 19521 1904
rect 19573 1852 19598 1904
rect 19494 1808 19598 1852
rect 17096 504 17364 526
rect 17096 388 17142 504
rect 17322 388 17364 504
rect 17096 356 17364 388
rect 17202 296 17304 356
rect 17206 -498 17286 296
rect 17090 -519 17396 -498
rect 17090 -575 17128 -519
rect 17184 -575 17208 -519
rect 17264 -575 17288 -519
rect 17344 -575 17396 -519
rect 17090 -594 17396 -575
rect 9712 -2000 9800 -1996
rect 16324 -1998 16416 -1704
rect 6312 -2002 6402 -2001
rect 16326 -2002 16416 -1998
rect 19697 -1999 19795 1906
rect 22840 2000 22946 2004
rect 26216 2165 26318 2202
rect 26216 2113 26240 2165
rect 26292 2113 26318 2165
rect 26216 2101 26318 2113
rect 26216 2049 26240 2101
rect 26292 2049 26318 2101
rect 26216 2037 26318 2049
rect 22840 1992 23096 2000
rect 22840 1940 22868 1992
rect 22920 1940 23096 1992
rect 22840 1928 23096 1940
rect 22840 1876 22868 1928
rect 22920 1904 23096 1928
rect 22920 1876 22946 1904
rect 22840 1864 22946 1876
rect 22840 1812 22868 1864
rect 22920 1812 22946 1864
rect 22840 1806 22946 1812
rect 20452 496 20718 524
rect 20452 380 20495 496
rect 20675 380 20718 496
rect 20452 346 20718 380
rect 20534 286 20636 346
rect 20549 -300 20627 286
rect 20436 -317 20742 -300
rect 20436 -373 20482 -317
rect 20538 -373 20562 -317
rect 20618 -373 20642 -317
rect 20698 -373 20742 -317
rect 20436 -396 20742 -373
rect 20549 -401 20627 -396
rect 23000 -2000 23096 1904
rect 26216 1985 26240 2037
rect 26292 2000 26318 2037
rect 26292 1985 26537 2000
rect 26216 1973 26537 1985
rect 26216 1921 26240 1973
rect 26292 1921 26537 1973
rect 26216 1910 26537 1921
rect 26216 1909 26318 1910
rect 26216 1857 26240 1909
rect 26292 1857 26318 1909
rect 26216 1812 26318 1857
rect 23824 509 24082 524
rect 23824 393 23861 509
rect 24041 393 24082 509
rect 23824 362 24082 393
rect 23898 -96 24000 362
rect 25858 249 26306 276
rect 25858 33 25893 249
rect 26269 33 26306 249
rect 25858 8 26306 33
rect 23800 -121 24106 -96
rect 23800 -177 23845 -121
rect 23901 -177 23925 -121
rect 23981 -177 24005 -121
rect 24061 -177 24106 -121
rect 23800 -202 24106 -177
rect 26447 -1698 26537 1910
rect 26446 -1996 26537 -1698
rect 26447 -1999 26537 -1996
<< via2 >>
rect -257 18 -41 154
rect 336 -1581 392 -1525
rect 416 -1581 472 -1525
rect 496 -1581 552 -1525
rect 3736 -1379 3792 -1323
rect 3816 -1379 3872 -1323
rect 3896 -1379 3952 -1323
rect 7056 -1179 7112 -1123
rect 7136 -1179 7192 -1123
rect 7216 -1179 7272 -1123
rect 10450 -975 10506 -919
rect 10530 -975 10586 -919
rect 10610 -975 10666 -919
rect 13740 -777 13796 -721
rect 13820 -777 13876 -721
rect 13900 -777 13956 -721
rect 17128 -575 17184 -519
rect 17208 -575 17264 -519
rect 17288 -575 17344 -519
rect 20482 -373 20538 -317
rect 20562 -373 20618 -317
rect 20642 -373 20698 -317
rect 25893 231 26269 249
rect 25893 51 25895 231
rect 25895 51 26267 231
rect 26267 51 26269 231
rect 25893 33 26269 51
rect 23845 -177 23901 -121
rect 23925 -177 23981 -121
rect 24005 -177 24061 -121
<< metal3 >>
rect -299 6684 1035 6802
rect 33400 4456 33702 4458
rect 27525 4396 33702 4456
rect 27525 3938 27585 4396
rect 30108 4264 33700 4324
rect 30108 4232 30169 4264
rect 30109 3924 30169 4232
rect 32828 4124 33704 4184
rect 32828 3996 32889 4124
rect 32829 3941 32889 3996
rect 23134 855 23454 910
rect -302 606 3320 730
rect 13144 614 13340 722
rect 23134 631 23176 855
rect 23400 631 23454 855
rect -300 602 -2 606
rect 23134 590 23454 631
rect 24366 606 24682 730
rect 25858 253 26306 276
rect -306 154 20 170
rect -306 18 -257 154
rect -41 18 20 154
rect -306 -4 20 18
rect 25858 29 25889 253
rect 26273 29 26306 253
rect 25858 8 26306 29
rect 26709 -96 26769 61
rect 23800 -117 24106 -96
rect 23800 -181 23841 -117
rect 23905 -181 23921 -117
rect 23985 -181 24001 -117
rect 24065 -181 24106 -117
rect 23800 -202 24106 -181
rect 26594 -118 26898 -96
rect 26594 -182 26634 -118
rect 26698 -182 26714 -118
rect 26778 -182 26794 -118
rect 26858 -182 26898 -118
rect 26594 -202 26898 -182
rect 27661 -300 27721 61
rect 20436 -313 20742 -300
rect 20436 -377 20478 -313
rect 20542 -377 20558 -313
rect 20622 -377 20638 -313
rect 20702 -377 20742 -313
rect 20436 -396 20742 -377
rect 27554 -314 27860 -300
rect 27554 -378 27599 -314
rect 27663 -378 27679 -314
rect 27743 -378 27759 -314
rect 27823 -378 27860 -314
rect 27554 -398 27860 -378
rect 17090 -515 17396 -498
rect 28613 -500 28673 68
rect 17090 -579 17124 -515
rect 17188 -579 17204 -515
rect 17268 -579 17284 -515
rect 17348 -579 17396 -515
rect 17090 -594 17396 -579
rect 28496 -518 28802 -500
rect 28496 -582 28531 -518
rect 28595 -582 28611 -518
rect 28675 -582 28691 -518
rect 28755 -582 28802 -518
rect 28496 -598 28802 -582
rect 13706 -717 14012 -698
rect 29701 -700 29761 61
rect 13706 -781 13736 -717
rect 13800 -781 13816 -717
rect 13880 -781 13896 -717
rect 13960 -781 14012 -717
rect 13706 -794 14012 -781
rect 29598 -713 29904 -700
rect 29598 -777 29637 -713
rect 29701 -777 29717 -713
rect 29781 -777 29797 -713
rect 29861 -777 29904 -713
rect 29598 -798 29904 -777
rect 29701 -800 29761 -798
rect 30653 -902 30713 61
rect 10406 -915 10712 -902
rect 10406 -979 10446 -915
rect 10510 -979 10526 -915
rect 10590 -979 10606 -915
rect 10670 -979 10712 -915
rect 10406 -998 10712 -979
rect 30546 -915 30852 -902
rect 30546 -979 30583 -915
rect 30647 -979 30663 -915
rect 30727 -979 30743 -915
rect 30807 -979 30852 -915
rect 30546 -1000 30852 -979
rect 30653 -1002 30713 -1000
rect 31605 -1098 31665 61
rect 7008 -1119 7314 -1100
rect 7008 -1183 7052 -1119
rect 7116 -1183 7132 -1119
rect 7196 -1183 7212 -1119
rect 7276 -1183 7314 -1119
rect 7008 -1196 7314 -1183
rect 31464 -1115 31770 -1098
rect 31464 -1179 31509 -1115
rect 31573 -1179 31589 -1115
rect 31653 -1179 31669 -1115
rect 31733 -1179 31770 -1115
rect 31464 -1196 31770 -1179
rect 31605 -1198 31665 -1196
rect 32693 -1300 32753 61
rect 3696 -1319 4002 -1300
rect 3696 -1383 3732 -1319
rect 3796 -1383 3812 -1319
rect 3876 -1383 3892 -1319
rect 3956 -1383 4002 -1319
rect 3696 -1396 4002 -1383
rect 32554 -1319 32860 -1300
rect 32554 -1383 32591 -1319
rect 32655 -1383 32671 -1319
rect 32735 -1383 32751 -1319
rect 32815 -1383 32860 -1319
rect 32554 -1398 32860 -1383
rect 32693 -1400 32753 -1398
rect 33445 -1502 33505 61
rect 298 -1521 604 -1504
rect 298 -1585 332 -1521
rect 396 -1585 412 -1521
rect 476 -1585 492 -1521
rect 556 -1585 604 -1521
rect 298 -1600 604 -1585
rect 33306 -1515 33612 -1502
rect 33306 -1579 33351 -1515
rect 33415 -1579 33431 -1515
rect 33495 -1579 33511 -1515
rect 33575 -1579 33612 -1515
rect 33306 -1600 33612 -1579
<< via3 >>
rect 23176 631 23400 855
rect 25889 249 26273 253
rect 25889 33 25893 249
rect 25893 33 26269 249
rect 26269 33 26273 249
rect 25889 29 26273 33
rect 23841 -121 23905 -117
rect 23841 -177 23845 -121
rect 23845 -177 23901 -121
rect 23901 -177 23905 -121
rect 23841 -181 23905 -177
rect 23921 -121 23985 -117
rect 23921 -177 23925 -121
rect 23925 -177 23981 -121
rect 23981 -177 23985 -121
rect 23921 -181 23985 -177
rect 24001 -121 24065 -117
rect 24001 -177 24005 -121
rect 24005 -177 24061 -121
rect 24061 -177 24065 -121
rect 24001 -181 24065 -177
rect 26634 -182 26698 -118
rect 26714 -182 26778 -118
rect 26794 -182 26858 -118
rect 20478 -317 20542 -313
rect 20478 -373 20482 -317
rect 20482 -373 20538 -317
rect 20538 -373 20542 -317
rect 20478 -377 20542 -373
rect 20558 -317 20622 -313
rect 20558 -373 20562 -317
rect 20562 -373 20618 -317
rect 20618 -373 20622 -317
rect 20558 -377 20622 -373
rect 20638 -317 20702 -313
rect 20638 -373 20642 -317
rect 20642 -373 20698 -317
rect 20698 -373 20702 -317
rect 20638 -377 20702 -373
rect 27599 -378 27663 -314
rect 27679 -378 27743 -314
rect 27759 -378 27823 -314
rect 17124 -519 17188 -515
rect 17124 -575 17128 -519
rect 17128 -575 17184 -519
rect 17184 -575 17188 -519
rect 17124 -579 17188 -575
rect 17204 -519 17268 -515
rect 17204 -575 17208 -519
rect 17208 -575 17264 -519
rect 17264 -575 17268 -519
rect 17204 -579 17268 -575
rect 17284 -519 17348 -515
rect 17284 -575 17288 -519
rect 17288 -575 17344 -519
rect 17344 -575 17348 -519
rect 17284 -579 17348 -575
rect 28531 -582 28595 -518
rect 28611 -582 28675 -518
rect 28691 -582 28755 -518
rect 13736 -721 13800 -717
rect 13736 -777 13740 -721
rect 13740 -777 13796 -721
rect 13796 -777 13800 -721
rect 13736 -781 13800 -777
rect 13816 -721 13880 -717
rect 13816 -777 13820 -721
rect 13820 -777 13876 -721
rect 13876 -777 13880 -721
rect 13816 -781 13880 -777
rect 13896 -721 13960 -717
rect 13896 -777 13900 -721
rect 13900 -777 13956 -721
rect 13956 -777 13960 -721
rect 13896 -781 13960 -777
rect 29637 -777 29701 -713
rect 29717 -777 29781 -713
rect 29797 -777 29861 -713
rect 10446 -919 10510 -915
rect 10446 -975 10450 -919
rect 10450 -975 10506 -919
rect 10506 -975 10510 -919
rect 10446 -979 10510 -975
rect 10526 -919 10590 -915
rect 10526 -975 10530 -919
rect 10530 -975 10586 -919
rect 10586 -975 10590 -919
rect 10526 -979 10590 -975
rect 10606 -919 10670 -915
rect 10606 -975 10610 -919
rect 10610 -975 10666 -919
rect 10666 -975 10670 -919
rect 10606 -979 10670 -975
rect 30583 -979 30647 -915
rect 30663 -979 30727 -915
rect 30743 -979 30807 -915
rect 7052 -1123 7116 -1119
rect 7052 -1179 7056 -1123
rect 7056 -1179 7112 -1123
rect 7112 -1179 7116 -1123
rect 7052 -1183 7116 -1179
rect 7132 -1123 7196 -1119
rect 7132 -1179 7136 -1123
rect 7136 -1179 7192 -1123
rect 7192 -1179 7196 -1123
rect 7132 -1183 7196 -1179
rect 7212 -1123 7276 -1119
rect 7212 -1179 7216 -1123
rect 7216 -1179 7272 -1123
rect 7272 -1179 7276 -1123
rect 7212 -1183 7276 -1179
rect 31509 -1179 31573 -1115
rect 31589 -1179 31653 -1115
rect 31669 -1179 31733 -1115
rect 3732 -1323 3796 -1319
rect 3732 -1379 3736 -1323
rect 3736 -1379 3792 -1323
rect 3792 -1379 3796 -1323
rect 3732 -1383 3796 -1379
rect 3812 -1323 3876 -1319
rect 3812 -1379 3816 -1323
rect 3816 -1379 3872 -1323
rect 3872 -1379 3876 -1323
rect 3812 -1383 3876 -1379
rect 3892 -1323 3956 -1319
rect 3892 -1379 3896 -1323
rect 3896 -1379 3952 -1323
rect 3952 -1379 3956 -1323
rect 3892 -1383 3956 -1379
rect 32591 -1383 32655 -1319
rect 32671 -1383 32735 -1319
rect 32751 -1383 32815 -1319
rect 332 -1525 396 -1521
rect 332 -1581 336 -1525
rect 336 -1581 392 -1525
rect 392 -1581 396 -1525
rect 332 -1585 396 -1581
rect 412 -1525 476 -1521
rect 412 -1581 416 -1525
rect 416 -1581 472 -1525
rect 472 -1581 476 -1525
rect 412 -1585 476 -1581
rect 492 -1525 556 -1521
rect 492 -1581 496 -1525
rect 496 -1581 552 -1525
rect 552 -1581 556 -1525
rect 492 -1585 556 -1581
rect 33351 -1579 33415 -1515
rect 33431 -1579 33495 -1515
rect 33511 -1579 33575 -1515
<< metal4 >>
rect 26562 3433 26798 3434
rect 23134 3113 26882 3433
rect 23134 855 23454 3113
rect 26562 3112 26798 3113
rect 26540 2793 26810 2798
rect 23134 631 23176 855
rect 23400 631 23454 855
rect 23134 592 23454 631
rect 26361 2474 26810 2793
rect 26361 273 26631 2474
rect 25855 253 26631 273
rect 25855 29 25889 253
rect 26273 29 26631 253
rect 25855 3 26631 29
rect -1 -117 33605 -100
rect -1 -181 23841 -117
rect 23905 -181 23921 -117
rect 23985 -181 24001 -117
rect 24065 -118 33605 -117
rect 24065 -181 26634 -118
rect -1 -182 26634 -181
rect 26698 -182 26714 -118
rect 26778 -182 26794 -118
rect 26858 -182 33605 -118
rect -1 -198 33605 -182
rect 0 -313 33606 -300
rect 0 -377 20478 -313
rect 20542 -377 20558 -313
rect 20622 -377 20638 -313
rect 20702 -314 33606 -313
rect 20702 -377 27599 -314
rect 0 -378 27599 -377
rect 27663 -378 27679 -314
rect 27743 -378 27759 -314
rect 27823 -378 33606 -314
rect 0 -398 33606 -378
rect 0 -515 33606 -500
rect 0 -579 17124 -515
rect 17188 -579 17204 -515
rect 17268 -579 17284 -515
rect 17348 -518 33606 -515
rect 17348 -579 28531 -518
rect 0 -582 28531 -579
rect 28595 -582 28611 -518
rect 28675 -582 28691 -518
rect 28755 -582 33606 -518
rect 0 -598 33606 -582
rect -2 -713 33604 -700
rect -2 -717 29637 -713
rect -2 -781 13736 -717
rect 13800 -781 13816 -717
rect 13880 -781 13896 -717
rect 13960 -777 29637 -717
rect 29701 -777 29717 -713
rect 29781 -777 29797 -713
rect 29861 -777 33604 -713
rect 13960 -781 33604 -777
rect -2 -798 33604 -781
rect 0 -915 33606 -902
rect 0 -979 10446 -915
rect 10510 -979 10526 -915
rect 10590 -979 10606 -915
rect 10670 -979 30583 -915
rect 30647 -979 30663 -915
rect 30727 -979 30743 -915
rect 30807 -979 33606 -915
rect 0 -1000 33606 -979
rect -2 -1115 33604 -1100
rect -2 -1119 31509 -1115
rect -2 -1183 7052 -1119
rect 7116 -1183 7132 -1119
rect 7196 -1183 7212 -1119
rect 7276 -1179 31509 -1119
rect 31573 -1179 31589 -1115
rect 31653 -1179 31669 -1115
rect 31733 -1179 33604 -1115
rect 7276 -1183 33604 -1179
rect -2 -1198 33604 -1183
rect 0 -1319 33606 -1300
rect 0 -1383 3732 -1319
rect 3796 -1383 3812 -1319
rect 3876 -1383 3892 -1319
rect 3956 -1383 32591 -1319
rect 32655 -1383 32671 -1319
rect 32735 -1383 32751 -1319
rect 32815 -1383 33606 -1319
rect 0 -1398 33606 -1383
rect 0 -1515 33606 -1502
rect 0 -1521 33351 -1515
rect 0 -1585 332 -1521
rect 396 -1585 412 -1521
rect 476 -1585 492 -1521
rect 556 -1579 33351 -1521
rect 33415 -1579 33431 -1515
rect 33495 -1579 33511 -1515
rect 33575 -1579 33606 -1515
rect 556 -1585 33606 -1579
rect 0 -1600 33606 -1585
use array_8ls_8tgwd_8sw  array_8ls_8tgwd_8sw_0
timestamp 1699926577
transform 1 0 13390 0 1 0
box -13390 -80 13065 11044
use decoder3to8  decoder3to8_0
timestamp 1699926577
transform 0 1 26261 -1 0 4030
box -274 394 4230 7249
<< labels >>
flabel metal2 s 26446 -1996 26536 -1698 0 FreeSans 1 0 0 0 VIN_0
port 1 nsew
flabel metal2 s 23004 -1998 23094 -1700 0 FreeSans 1 0 0 0 VIN_1
port 2 nsew
flabel metal2 s 19698 -1998 19788 -1700 0 FreeSans 1 0 0 0 VIN_2
port 3 nsew
flabel metal2 s 16326 -2002 16416 -1704 0 FreeSans 1 0 0 0 VIN_3
port 4 nsew
flabel metal2 s 13012 -1996 13102 -1698 0 FreeSans 1 0 0 0 VIN_4
port 5 nsew
flabel metal2 s 9712 -1996 9802 -1698 0 FreeSans 1 0 0 0 VIN_5
port 6 nsew
flabel metal2 s 6312 -2002 6402 -1704 0 FreeSans 1 0 0 0 VIN_6
port 7 nsew
flabel metal2 s 2908 -2006 2998 -1708 0 FreeSans 1 0 0 0 VIN_7
port 8 nsew
flabel metal3 s -300 602 -2 730 0 FreeSans 1 0 0 0 DVDD
port 9 nsew
flabel metal3 s 13144 614 13340 722 0 FreeSans 1 0 0 0 DVDD
port 9 nsew
flabel metal3 s 33396 4124 33704 4184 0 FreeSans 1 0 0 0 B0
port 10 nsew
flabel metal3 s 33398 4266 33700 4324 0 FreeSans 1 0 0 0 B1
port 11 nsew
flabel metal3 s 33400 4400 33702 4458 0 FreeSans 1 0 0 0 B2
port 12 nsew
flabel metal3 s -306 -4 20 170 0 FreeSans 1 0 0 0 DVSS
port 13 nsew
flabel metal3 s -298 6686 2 6800 0 FreeSans 1 0 0 0 VDD
port 14 nsew
flabel metal2 s 12900 10934 13304 11042 0 FreeSans 49 0 0 0 VO
port 15 nsew
<< end >>
