magic
tech sky130A
magscale 1 2
timestamp 1699926577
<< pwell >>
rect -418 -748 418 748
<< mvnmos >>
rect -200 -500 200 500
<< mvndiff >>
rect -258 459 -200 500
rect -258 425 -246 459
rect -212 425 -200 459
rect -258 391 -200 425
rect -258 357 -246 391
rect -212 357 -200 391
rect -258 323 -200 357
rect -258 289 -246 323
rect -212 289 -200 323
rect -258 255 -200 289
rect -258 221 -246 255
rect -212 221 -200 255
rect -258 187 -200 221
rect -258 153 -246 187
rect -212 153 -200 187
rect -258 119 -200 153
rect -258 85 -246 119
rect -212 85 -200 119
rect -258 51 -200 85
rect -258 17 -246 51
rect -212 17 -200 51
rect -258 -17 -200 17
rect -258 -51 -246 -17
rect -212 -51 -200 -17
rect -258 -85 -200 -51
rect -258 -119 -246 -85
rect -212 -119 -200 -85
rect -258 -153 -200 -119
rect -258 -187 -246 -153
rect -212 -187 -200 -153
rect -258 -221 -200 -187
rect -258 -255 -246 -221
rect -212 -255 -200 -221
rect -258 -289 -200 -255
rect -258 -323 -246 -289
rect -212 -323 -200 -289
rect -258 -357 -200 -323
rect -258 -391 -246 -357
rect -212 -391 -200 -357
rect -258 -425 -200 -391
rect -258 -459 -246 -425
rect -212 -459 -200 -425
rect -258 -500 -200 -459
rect 200 459 258 500
rect 200 425 212 459
rect 246 425 258 459
rect 200 391 258 425
rect 200 357 212 391
rect 246 357 258 391
rect 200 323 258 357
rect 200 289 212 323
rect 246 289 258 323
rect 200 255 258 289
rect 200 221 212 255
rect 246 221 258 255
rect 200 187 258 221
rect 200 153 212 187
rect 246 153 258 187
rect 200 119 258 153
rect 200 85 212 119
rect 246 85 258 119
rect 200 51 258 85
rect 200 17 212 51
rect 246 17 258 51
rect 200 -17 258 17
rect 200 -51 212 -17
rect 246 -51 258 -17
rect 200 -85 258 -51
rect 200 -119 212 -85
rect 246 -119 258 -85
rect 200 -153 258 -119
rect 200 -187 212 -153
rect 246 -187 258 -153
rect 200 -221 258 -187
rect 200 -255 212 -221
rect 246 -255 258 -221
rect 200 -289 258 -255
rect 200 -323 212 -289
rect 246 -323 258 -289
rect 200 -357 258 -323
rect 200 -391 212 -357
rect 246 -391 258 -357
rect 200 -425 258 -391
rect 200 -459 212 -425
rect 246 -459 258 -425
rect 200 -500 258 -459
<< mvndiffc >>
rect -246 425 -212 459
rect -246 357 -212 391
rect -246 289 -212 323
rect -246 221 -212 255
rect -246 153 -212 187
rect -246 85 -212 119
rect -246 17 -212 51
rect -246 -51 -212 -17
rect -246 -119 -212 -85
rect -246 -187 -212 -153
rect -246 -255 -212 -221
rect -246 -323 -212 -289
rect -246 -391 -212 -357
rect -246 -459 -212 -425
rect 212 425 246 459
rect 212 357 246 391
rect 212 289 246 323
rect 212 221 246 255
rect 212 153 246 187
rect 212 85 246 119
rect 212 17 246 51
rect 212 -51 246 -17
rect 212 -119 246 -85
rect 212 -187 246 -153
rect 212 -255 246 -221
rect 212 -323 246 -289
rect 212 -391 246 -357
rect 212 -459 246 -425
<< mvpsubdiff >>
rect -392 710 392 722
rect -392 676 -255 710
rect -221 676 -187 710
rect -153 676 -119 710
rect -85 676 -51 710
rect -17 676 17 710
rect 51 676 85 710
rect 119 676 153 710
rect 187 676 221 710
rect 255 676 392 710
rect -392 664 392 676
rect -392 595 -334 664
rect -392 561 -380 595
rect -346 561 -334 595
rect 334 595 392 664
rect -392 527 -334 561
rect -392 493 -380 527
rect -346 493 -334 527
rect 334 561 346 595
rect 380 561 392 595
rect 334 527 392 561
rect -392 459 -334 493
rect -392 425 -380 459
rect -346 425 -334 459
rect -392 391 -334 425
rect -392 357 -380 391
rect -346 357 -334 391
rect -392 323 -334 357
rect -392 289 -380 323
rect -346 289 -334 323
rect -392 255 -334 289
rect -392 221 -380 255
rect -346 221 -334 255
rect -392 187 -334 221
rect -392 153 -380 187
rect -346 153 -334 187
rect -392 119 -334 153
rect -392 85 -380 119
rect -346 85 -334 119
rect -392 51 -334 85
rect -392 17 -380 51
rect -346 17 -334 51
rect -392 -17 -334 17
rect -392 -51 -380 -17
rect -346 -51 -334 -17
rect -392 -85 -334 -51
rect -392 -119 -380 -85
rect -346 -119 -334 -85
rect -392 -153 -334 -119
rect -392 -187 -380 -153
rect -346 -187 -334 -153
rect -392 -221 -334 -187
rect -392 -255 -380 -221
rect -346 -255 -334 -221
rect -392 -289 -334 -255
rect -392 -323 -380 -289
rect -346 -323 -334 -289
rect -392 -357 -334 -323
rect -392 -391 -380 -357
rect -346 -391 -334 -357
rect -392 -425 -334 -391
rect -392 -459 -380 -425
rect -346 -459 -334 -425
rect -392 -493 -334 -459
rect -392 -527 -380 -493
rect -346 -527 -334 -493
rect 334 493 346 527
rect 380 493 392 527
rect 334 459 392 493
rect 334 425 346 459
rect 380 425 392 459
rect 334 391 392 425
rect 334 357 346 391
rect 380 357 392 391
rect 334 323 392 357
rect 334 289 346 323
rect 380 289 392 323
rect 334 255 392 289
rect 334 221 346 255
rect 380 221 392 255
rect 334 187 392 221
rect 334 153 346 187
rect 380 153 392 187
rect 334 119 392 153
rect 334 85 346 119
rect 380 85 392 119
rect 334 51 392 85
rect 334 17 346 51
rect 380 17 392 51
rect 334 -17 392 17
rect 334 -51 346 -17
rect 380 -51 392 -17
rect 334 -85 392 -51
rect 334 -119 346 -85
rect 380 -119 392 -85
rect 334 -153 392 -119
rect 334 -187 346 -153
rect 380 -187 392 -153
rect 334 -221 392 -187
rect 334 -255 346 -221
rect 380 -255 392 -221
rect 334 -289 392 -255
rect 334 -323 346 -289
rect 380 -323 392 -289
rect 334 -357 392 -323
rect 334 -391 346 -357
rect 380 -391 392 -357
rect 334 -425 392 -391
rect 334 -459 346 -425
rect 380 -459 392 -425
rect 334 -493 392 -459
rect -392 -561 -334 -527
rect -392 -595 -380 -561
rect -346 -595 -334 -561
rect 334 -527 346 -493
rect 380 -527 392 -493
rect 334 -561 392 -527
rect -392 -664 -334 -595
rect 334 -595 346 -561
rect 380 -595 392 -561
rect 334 -664 392 -595
rect -392 -676 392 -664
rect -392 -710 -255 -676
rect -221 -710 -187 -676
rect -153 -710 -119 -676
rect -85 -710 -51 -676
rect -17 -710 17 -676
rect 51 -710 85 -676
rect 119 -710 153 -676
rect 187 -710 221 -676
rect 255 -710 392 -676
rect -392 -722 392 -710
<< mvpsubdiffcont >>
rect -255 676 -221 710
rect -187 676 -153 710
rect -119 676 -85 710
rect -51 676 -17 710
rect 17 676 51 710
rect 85 676 119 710
rect 153 676 187 710
rect 221 676 255 710
rect -380 561 -346 595
rect -380 493 -346 527
rect 346 561 380 595
rect -380 425 -346 459
rect -380 357 -346 391
rect -380 289 -346 323
rect -380 221 -346 255
rect -380 153 -346 187
rect -380 85 -346 119
rect -380 17 -346 51
rect -380 -51 -346 -17
rect -380 -119 -346 -85
rect -380 -187 -346 -153
rect -380 -255 -346 -221
rect -380 -323 -346 -289
rect -380 -391 -346 -357
rect -380 -459 -346 -425
rect -380 -527 -346 -493
rect 346 493 380 527
rect 346 425 380 459
rect 346 357 380 391
rect 346 289 380 323
rect 346 221 380 255
rect 346 153 380 187
rect 346 85 380 119
rect 346 17 380 51
rect 346 -51 380 -17
rect 346 -119 380 -85
rect 346 -187 380 -153
rect 346 -255 380 -221
rect 346 -323 380 -289
rect 346 -391 380 -357
rect 346 -459 380 -425
rect -380 -595 -346 -561
rect 346 -527 380 -493
rect 346 -595 380 -561
rect -255 -710 -221 -676
rect -187 -710 -153 -676
rect -119 -710 -85 -676
rect -51 -710 -17 -676
rect 17 -710 51 -676
rect 85 -710 119 -676
rect 153 -710 187 -676
rect 221 -710 255 -676
<< poly >>
rect -200 572 200 588
rect -200 538 -153 572
rect -119 538 -85 572
rect -51 538 -17 572
rect 17 538 51 572
rect 85 538 119 572
rect 153 538 200 572
rect -200 500 200 538
rect -200 -538 200 -500
rect -200 -572 -153 -538
rect -119 -572 -85 -538
rect -51 -572 -17 -538
rect 17 -572 51 -538
rect 85 -572 119 -538
rect 153 -572 200 -538
rect -200 -588 200 -572
<< polycont >>
rect -153 538 -119 572
rect -85 538 -51 572
rect -17 538 17 572
rect 51 538 85 572
rect 119 538 153 572
rect -153 -572 -119 -538
rect -85 -572 -51 -538
rect -17 -572 17 -538
rect 51 -572 85 -538
rect 119 -572 153 -538
<< locali >>
rect -380 676 -255 710
rect -221 676 -187 710
rect -153 676 -119 710
rect -85 676 -51 710
rect -17 676 17 710
rect 51 676 85 710
rect 119 676 153 710
rect 187 676 221 710
rect 255 676 380 710
rect -380 595 -346 676
rect 346 665 380 676
rect 346 595 380 631
rect -380 527 -346 561
rect -200 538 -161 572
rect -119 538 -89 572
rect -51 538 -17 572
rect 17 538 51 572
rect 89 538 119 572
rect 161 538 200 572
rect 346 527 380 559
rect -380 459 -346 493
rect -380 391 -346 425
rect -380 323 -346 357
rect -380 255 -346 289
rect -380 187 -346 221
rect -380 119 -346 153
rect -380 51 -346 85
rect -380 -17 -346 17
rect -380 -85 -346 -51
rect -380 -153 -346 -119
rect -380 -221 -346 -187
rect -380 -289 -346 -255
rect -380 -357 -346 -323
rect -380 -425 -346 -391
rect -380 -493 -346 -459
rect -246 485 -212 504
rect -246 413 -212 425
rect -246 341 -212 357
rect -246 269 -212 289
rect -246 197 -212 221
rect -246 125 -212 153
rect -246 53 -212 85
rect -246 -17 -212 17
rect -246 -85 -212 -53
rect -246 -153 -212 -125
rect -246 -221 -212 -197
rect -246 -289 -212 -269
rect -246 -357 -212 -341
rect -246 -425 -212 -413
rect -246 -504 -212 -485
rect 212 485 246 504
rect 212 413 246 425
rect 212 341 246 357
rect 212 269 246 289
rect 212 197 246 221
rect 212 125 246 153
rect 212 53 246 85
rect 212 -17 246 17
rect 212 -85 246 -53
rect 212 -153 246 -125
rect 212 -221 246 -197
rect 212 -289 246 -269
rect 212 -357 246 -341
rect 212 -425 246 -413
rect 212 -504 246 -485
rect 346 459 380 487
rect 346 391 380 415
rect 346 323 380 343
rect 346 255 380 271
rect 346 187 380 199
rect 346 119 380 127
rect 346 51 380 55
rect 346 -55 380 -51
rect 346 -127 380 -119
rect 346 -199 380 -187
rect 346 -271 380 -255
rect 346 -343 380 -323
rect 346 -415 380 -391
rect 346 -487 380 -459
rect -380 -561 -346 -527
rect -200 -572 -161 -538
rect -119 -572 -89 -538
rect -51 -572 -17 -538
rect 17 -572 51 -538
rect 89 -572 119 -538
rect 161 -572 200 -538
rect 346 -559 380 -527
rect -380 -676 -346 -595
rect 346 -631 380 -595
rect 346 -676 380 -665
rect -380 -710 -255 -676
rect -221 -710 -187 -676
rect -153 -710 -119 -676
rect -85 -710 -51 -676
rect -17 -710 17 -676
rect 51 -710 85 -676
rect 119 -710 153 -676
rect 187 -710 221 -676
rect 255 -710 380 -676
<< viali >>
rect 346 631 380 665
rect -161 538 -153 572
rect -153 538 -127 572
rect -89 538 -85 572
rect -85 538 -55 572
rect -17 538 17 572
rect 55 538 85 572
rect 85 538 89 572
rect 127 538 153 572
rect 153 538 161 572
rect 346 561 380 593
rect 346 559 380 561
rect -246 459 -212 485
rect -246 451 -212 459
rect -246 391 -212 413
rect -246 379 -212 391
rect -246 323 -212 341
rect -246 307 -212 323
rect -246 255 -212 269
rect -246 235 -212 255
rect -246 187 -212 197
rect -246 163 -212 187
rect -246 119 -212 125
rect -246 91 -212 119
rect -246 51 -212 53
rect -246 19 -212 51
rect -246 -51 -212 -19
rect -246 -53 -212 -51
rect -246 -119 -212 -91
rect -246 -125 -212 -119
rect -246 -187 -212 -163
rect -246 -197 -212 -187
rect -246 -255 -212 -235
rect -246 -269 -212 -255
rect -246 -323 -212 -307
rect -246 -341 -212 -323
rect -246 -391 -212 -379
rect -246 -413 -212 -391
rect -246 -459 -212 -451
rect -246 -485 -212 -459
rect 212 459 246 485
rect 212 451 246 459
rect 212 391 246 413
rect 212 379 246 391
rect 212 323 246 341
rect 212 307 246 323
rect 212 255 246 269
rect 212 235 246 255
rect 212 187 246 197
rect 212 163 246 187
rect 212 119 246 125
rect 212 91 246 119
rect 212 51 246 53
rect 212 19 246 51
rect 212 -51 246 -19
rect 212 -53 246 -51
rect 212 -119 246 -91
rect 212 -125 246 -119
rect 212 -187 246 -163
rect 212 -197 246 -187
rect 212 -255 246 -235
rect 212 -269 246 -255
rect 212 -323 246 -307
rect 212 -341 246 -323
rect 212 -391 246 -379
rect 212 -413 246 -391
rect 212 -459 246 -451
rect 212 -485 246 -459
rect 346 493 380 521
rect 346 487 380 493
rect 346 425 380 449
rect 346 415 380 425
rect 346 357 380 377
rect 346 343 380 357
rect 346 289 380 305
rect 346 271 380 289
rect 346 221 380 233
rect 346 199 380 221
rect 346 153 380 161
rect 346 127 380 153
rect 346 85 380 89
rect 346 55 380 85
rect 346 -17 380 17
rect 346 -85 380 -55
rect 346 -89 380 -85
rect 346 -153 380 -127
rect 346 -161 380 -153
rect 346 -221 380 -199
rect 346 -233 380 -221
rect 346 -289 380 -271
rect 346 -305 380 -289
rect 346 -357 380 -343
rect 346 -377 380 -357
rect 346 -425 380 -415
rect 346 -449 380 -425
rect 346 -493 380 -487
rect 346 -521 380 -493
rect -161 -572 -153 -538
rect -153 -572 -127 -538
rect -89 -572 -85 -538
rect -85 -572 -55 -538
rect -17 -572 17 -538
rect 55 -572 85 -538
rect 85 -572 89 -538
rect 127 -572 153 -538
rect 153 -572 161 -538
rect 346 -561 380 -559
rect 346 -593 380 -561
rect 346 -665 380 -631
<< metal1 >>
rect 340 665 386 688
rect 340 631 346 665
rect 380 631 386 665
rect 340 593 386 631
rect -196 572 196 578
rect -196 538 -161 572
rect -127 538 -89 572
rect -55 538 -17 572
rect 17 538 55 572
rect 89 538 127 572
rect 161 538 196 572
rect -196 532 196 538
rect 340 559 346 593
rect 380 559 386 593
rect 340 521 386 559
rect -252 485 -206 500
rect -252 451 -246 485
rect -212 451 -206 485
rect -252 413 -206 451
rect -252 379 -246 413
rect -212 379 -206 413
rect -252 341 -206 379
rect -252 307 -246 341
rect -212 307 -206 341
rect -252 269 -206 307
rect -252 235 -246 269
rect -212 235 -206 269
rect -252 197 -206 235
rect -252 163 -246 197
rect -212 163 -206 197
rect -252 125 -206 163
rect -252 91 -246 125
rect -212 91 -206 125
rect -252 53 -206 91
rect -252 19 -246 53
rect -212 19 -206 53
rect -252 -19 -206 19
rect -252 -53 -246 -19
rect -212 -53 -206 -19
rect -252 -91 -206 -53
rect -252 -125 -246 -91
rect -212 -125 -206 -91
rect -252 -163 -206 -125
rect -252 -197 -246 -163
rect -212 -197 -206 -163
rect -252 -235 -206 -197
rect -252 -269 -246 -235
rect -212 -269 -206 -235
rect -252 -307 -206 -269
rect -252 -341 -246 -307
rect -212 -341 -206 -307
rect -252 -379 -206 -341
rect -252 -413 -246 -379
rect -212 -413 -206 -379
rect -252 -451 -206 -413
rect -252 -485 -246 -451
rect -212 -485 -206 -451
rect -252 -500 -206 -485
rect 206 485 252 500
rect 206 451 212 485
rect 246 451 252 485
rect 206 413 252 451
rect 206 379 212 413
rect 246 379 252 413
rect 206 341 252 379
rect 206 307 212 341
rect 246 307 252 341
rect 206 269 252 307
rect 206 235 212 269
rect 246 235 252 269
rect 206 197 252 235
rect 206 163 212 197
rect 246 163 252 197
rect 206 125 252 163
rect 206 91 212 125
rect 246 91 252 125
rect 206 53 252 91
rect 206 19 212 53
rect 246 19 252 53
rect 206 -19 252 19
rect 206 -53 212 -19
rect 246 -53 252 -19
rect 206 -91 252 -53
rect 206 -125 212 -91
rect 246 -125 252 -91
rect 206 -163 252 -125
rect 206 -197 212 -163
rect 246 -197 252 -163
rect 206 -235 252 -197
rect 206 -269 212 -235
rect 246 -269 252 -235
rect 206 -307 252 -269
rect 206 -341 212 -307
rect 246 -341 252 -307
rect 206 -379 252 -341
rect 206 -413 212 -379
rect 246 -413 252 -379
rect 206 -451 252 -413
rect 206 -485 212 -451
rect 246 -485 252 -451
rect 206 -500 252 -485
rect 340 487 346 521
rect 380 487 386 521
rect 340 449 386 487
rect 340 415 346 449
rect 380 415 386 449
rect 340 377 386 415
rect 340 343 346 377
rect 380 343 386 377
rect 340 305 386 343
rect 340 271 346 305
rect 380 271 386 305
rect 340 233 386 271
rect 340 199 346 233
rect 380 199 386 233
rect 340 161 386 199
rect 340 127 346 161
rect 380 127 386 161
rect 340 89 386 127
rect 340 55 346 89
rect 380 55 386 89
rect 340 17 386 55
rect 340 -17 346 17
rect 380 -17 386 17
rect 340 -55 386 -17
rect 340 -89 346 -55
rect 380 -89 386 -55
rect 340 -127 386 -89
rect 340 -161 346 -127
rect 380 -161 386 -127
rect 340 -199 386 -161
rect 340 -233 346 -199
rect 380 -233 386 -199
rect 340 -271 386 -233
rect 340 -305 346 -271
rect 380 -305 386 -271
rect 340 -343 386 -305
rect 340 -377 346 -343
rect 380 -377 386 -343
rect 340 -415 386 -377
rect 340 -449 346 -415
rect 380 -449 386 -415
rect 340 -487 386 -449
rect 340 -521 346 -487
rect 380 -521 386 -487
rect -196 -538 196 -532
rect -196 -572 -161 -538
rect -127 -572 -89 -538
rect -55 -572 -17 -538
rect 17 -572 55 -538
rect 89 -572 127 -538
rect 161 -572 196 -538
rect -196 -578 196 -572
rect 340 -559 386 -521
rect 340 -593 346 -559
rect 380 -593 386 -559
rect 340 -631 386 -593
rect 340 -665 346 -631
rect 380 -665 386 -631
rect 340 -688 386 -665
<< properties >>
string FIXED_BBOX -363 -693 363 693
<< end >>
