VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO EF_ADCS1008NC
  CLASS BLOCK ;
  FOREIGN EF_ADCS1008NC ;
  ORIGIN -28.140 -1837.465 ;
  SIZE 348.430 BY 531.590 ;
  PIN B[0]
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 207.260 2338.105 208.800 2338.405 ;
    END
  END B[0]
  PIN B[1]
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 207.250 2337.415 208.790 2337.715 ;
    END
  END B[1]
  PIN B[2]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 207.270 2336.745 208.810 2337.045 ;
    END
  END B[2]
  PIN VIN[0]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 172.510 2367.515 172.965 2369.005 ;
    END
  END VIN[0]
  PIN VIN[1]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 155.290 2367.515 155.770 2369.025 ;
    END
  END VIN[1]
  PIN VIN[2]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 138.770 2367.535 139.250 2369.045 ;
    END
  END VIN[2]
  PIN VIN[3]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 121.890 2367.555 122.350 2369.035 ;
    END
  END VIN[3]
  PIN VIN[4]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 105.340 2367.525 105.800 2369.005 ;
    END
  END VIN[4]
  PIN VIN[5]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 88.820 2367.535 89.280 2369.015 ;
    END
  END VIN[5]
  PIN VIN[6]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 71.830 2367.535 72.290 2369.015 ;
    END
  END VIN[6]
  PIN VIN[7]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 54.840 2367.555 55.300 2369.035 ;
    END
  END VIN[7]
  PIN HOLD
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.360000 ;
    PORT
      LAYER met1 ;
        RECT 38.570 2285.280 39.570 2286.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.710 2285.295 35.860 2286.305 ;
    END
  END HOLD
  PIN CMP
    ANTENNADIFFAREA 0.492900 ;
    PORT
      LAYER met3 ;
        RECT 206.690 2261.575 208.760 2262.565 ;
    END
  END CMP
  PIN DATA[9]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 38.720 2171.045 44.480 2171.925 ;
    END
  END DATA[9]
  PIN DATA[8]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 38.740 2137.415 44.500 2138.295 ;
    END
  END DATA[8]
  PIN DATA[7]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 38.700 2103.835 44.460 2104.715 ;
    END
  END DATA[7]
  PIN DATA[6]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 38.760 2070.365 44.520 2071.245 ;
    END
  END DATA[6]
  PIN DATA[5]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 38.780 2036.515 44.540 2037.395 ;
    END
  END DATA[5]
  PIN DATA[0]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 38.720 2001.585 44.480 2002.465 ;
    END
  END DATA[0]
  PIN DATA[1]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 38.760 1968.055 44.520 1968.935 ;
    END
  END DATA[1]
  PIN DATA[2]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 38.740 1934.455 44.500 1935.335 ;
    END
  END DATA[2]
  PIN DATA[3]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 38.700 1900.945 44.460 1901.825 ;
    END
  END DATA[3]
  PIN DATA[4]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 38.720 1867.055 44.480 1867.935 ;
    END
  END DATA[4]
  PIN VH
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met3 ;
        RECT 38.720 2031.955 44.480 2032.835 ;
    END
  END VH
  PIN VL
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met3 ;
        RECT 38.670 2029.625 44.430 2030.505 ;
    END
  END VL
  PIN RST
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER met3 ;
        RECT 36.720 2228.595 40.820 2229.605 ;
    END
  END RST
  PIN DVDD
    ANTENNAGATEAREA 47.261497 ;
    ANTENNADIFFAREA 93.596451 ;
    PORT
      LAYER met3 ;
        RECT 38.760 1859.355 45.950 1861.345 ;
    END
  END DVDD
  PIN DVSS
    ANTENNAGATEAREA 74.759102 ;
    ANTENNADIFFAREA 1023.766663 ;
    PORT
      LAYER met3 ;
        RECT 38.730 1856.685 45.920 1858.675 ;
    END
  END DVSS
  PIN VSS
    ANTENNAGATEAREA 130.500000 ;
    ANTENNADIFFAREA 621.362671 ;
    PORT
      LAYER met3 ;
        RECT 38.720 1851.465 46.130 1853.365 ;
    END
  END VSS
  PIN VDD
    ANTENNAGATEAREA 100.000000 ;
    ANTENNADIFFAREA 2509.495605 ;
    PORT
      LAYER met3 ;
        RECT 38.840 1854.225 46.140 1856.165 ;
    END
  END VDD
  PIN EN
    ANTENNAGATEAREA 1.752000 ;
    ANTENNADIFFAREA 1.080000 ;
    PORT
      LAYER met3 ;
        RECT 32.710 2264.065 35.500 2264.995 ;
    END
  END EN
  OBS
      LAYER li1 ;
        RECT 39.935 1865.505 280.620 2358.820 ;
      LAYER met1 ;
        RECT 32.755 2286.560 281.315 2359.025 ;
        RECT 32.755 2285.000 38.290 2286.560 ;
        RECT 39.850 2285.000 281.315 2286.560 ;
        RECT 32.755 1863.190 281.315 2285.000 ;
      LAYER met2 ;
        RECT 32.710 2367.275 54.560 2369.055 ;
        RECT 55.580 2367.275 71.550 2369.055 ;
        RECT 32.710 2367.255 71.550 2367.275 ;
        RECT 72.570 2367.255 88.540 2369.055 ;
        RECT 89.560 2367.255 105.060 2369.055 ;
        RECT 32.710 2367.245 105.060 2367.255 ;
        RECT 106.080 2367.275 121.610 2369.055 ;
        RECT 122.630 2367.275 138.490 2369.055 ;
        RECT 106.080 2367.255 138.490 2367.275 ;
        RECT 139.530 2367.255 155.010 2369.055 ;
        RECT 106.080 2367.245 155.010 2367.255 ;
        RECT 32.710 2367.235 155.010 2367.245 ;
        RECT 156.050 2367.235 172.230 2369.055 ;
        RECT 173.245 2367.235 279.000 2369.055 ;
        RECT 32.710 1863.190 279.000 2367.235 ;
      LAYER met3 ;
        RECT 32.700 2338.805 376.570 2367.025 ;
        RECT 32.700 2338.115 206.860 2338.805 ;
        RECT 32.700 2337.015 206.850 2338.115 ;
        RECT 209.200 2337.705 376.570 2338.805 ;
        RECT 209.190 2337.445 376.570 2337.705 ;
        RECT 32.700 2336.345 206.870 2337.015 ;
        RECT 209.210 2336.345 376.570 2337.445 ;
        RECT 32.700 2286.705 376.570 2336.345 ;
        RECT 36.260 2284.895 376.570 2286.705 ;
        RECT 32.700 2265.395 376.570 2284.895 ;
        RECT 35.900 2263.665 376.570 2265.395 ;
        RECT 32.700 2262.965 376.570 2263.665 ;
        RECT 32.700 2261.175 206.290 2262.965 ;
        RECT 209.160 2261.175 376.570 2262.965 ;
        RECT 32.700 2230.005 376.570 2261.175 ;
        RECT 32.700 2228.195 36.320 2230.005 ;
        RECT 41.220 2228.195 376.570 2230.005 ;
        RECT 32.700 2172.325 376.570 2228.195 ;
        RECT 32.700 2170.645 38.320 2172.325 ;
        RECT 44.880 2170.645 376.570 2172.325 ;
        RECT 32.700 2138.695 376.570 2170.645 ;
        RECT 32.700 2137.015 38.340 2138.695 ;
        RECT 44.900 2137.015 376.570 2138.695 ;
        RECT 32.700 2105.115 376.570 2137.015 ;
        RECT 32.700 2103.435 38.300 2105.115 ;
        RECT 44.860 2103.435 376.570 2105.115 ;
        RECT 32.700 2071.645 376.570 2103.435 ;
        RECT 32.700 2069.965 38.360 2071.645 ;
        RECT 44.920 2069.965 376.570 2071.645 ;
        RECT 32.700 2037.795 376.570 2069.965 ;
        RECT 32.700 2036.115 38.380 2037.795 ;
        RECT 44.940 2036.115 376.570 2037.795 ;
        RECT 32.700 2033.235 376.570 2036.115 ;
        RECT 32.700 2031.555 38.320 2033.235 ;
        RECT 44.880 2031.555 376.570 2033.235 ;
        RECT 32.700 2030.905 376.570 2031.555 ;
        RECT 32.700 2029.225 38.270 2030.905 ;
        RECT 44.830 2029.225 376.570 2030.905 ;
        RECT 32.700 2002.865 376.570 2029.225 ;
        RECT 32.700 2001.185 38.320 2002.865 ;
        RECT 44.880 2001.185 376.570 2002.865 ;
        RECT 32.700 1969.335 376.570 2001.185 ;
        RECT 32.700 1967.655 38.360 1969.335 ;
        RECT 44.920 1967.655 376.570 1969.335 ;
        RECT 32.700 1935.735 376.570 1967.655 ;
        RECT 32.700 1934.055 38.340 1935.735 ;
        RECT 44.900 1934.055 376.570 1935.735 ;
        RECT 32.700 1902.225 376.570 1934.055 ;
        RECT 32.700 1900.545 38.300 1902.225 ;
        RECT 44.860 1900.545 376.570 1902.225 ;
        RECT 32.700 1868.335 376.570 1900.545 ;
        RECT 32.700 1866.655 38.320 1868.335 ;
        RECT 44.880 1866.655 376.570 1868.335 ;
        RECT 32.700 1861.745 376.570 1866.655 ;
        RECT 32.700 1859.075 38.360 1861.745 ;
        RECT 32.700 1856.285 38.330 1859.075 ;
        RECT 46.350 1858.955 376.570 1861.745 ;
        RECT 46.320 1856.565 376.570 1858.955 ;
        RECT 32.700 1853.825 38.440 1856.285 ;
        RECT 46.540 1853.825 376.570 1856.565 ;
        RECT 32.700 1853.765 376.570 1853.825 ;
        RECT 32.700 1851.430 38.320 1853.765 ;
        RECT 46.530 1851.430 376.570 1853.765 ;
      LAYER met4 ;
        RECT 36.580 1851.430 376.400 2367.025 ;
      LAYER met5 ;
        RECT 49.645 2235.910 203.675 2358.340 ;
  END
END EF_ADCS1008NC
END LIBRARY

