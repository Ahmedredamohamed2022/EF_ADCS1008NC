magic
tech sky130A
magscale 1 2
timestamp 1699926577
<< metal3 >>
rect 2013 -17007 3394 -16918
rect 4122 -17007 6780 -16918
rect 7508 -17007 10166 -16918
rect 10894 -17007 13552 -16918
rect 14280 -17007 16938 -16918
rect 17666 -17007 19047 -16918
rect 2013 -18296 3394 -18207
rect 4122 -18296 6780 -18207
rect 7508 -18296 10166 -18207
rect 10894 -18296 13552 -18207
rect 14280 -18296 16938 -18207
rect 17666 -18296 19047 -18207
rect 2013 -19585 3394 -19496
rect 4122 -19585 6780 -19496
rect 7508 -19585 10166 -19496
rect 10894 -19585 13552 -19496
rect 14280 -19585 16938 -19496
rect 17666 -19585 19047 -19496
rect 2013 -20874 3394 -20785
rect 4122 -20874 6780 -20785
rect 7508 -20874 10166 -20785
rect 10894 -20874 13552 -20785
rect 14280 -20874 16938 -20785
rect 17666 -20874 19047 -20785
rect 2013 -22163 3394 -22074
rect 4122 -22163 6780 -22074
rect 7508 -22163 10166 -22074
rect 10894 -22163 13552 -22074
rect 14280 -22163 16938 -22074
rect 17666 -22163 19047 -22074
rect 2013 -23452 3395 -23363
rect 4122 -23452 6780 -23363
rect 7508 -23452 10166 -23363
rect 10894 -23452 13552 -23363
rect 14280 -23452 16938 -23363
rect 17666 -23452 19047 -23363
rect 2013 -24741 3394 -24652
rect 4122 -24741 6780 -24652
rect 7508 -24741 10166 -24652
rect 10894 -24741 13552 -24652
rect 14280 -24741 16938 -24652
rect 17666 -24741 19047 -24652
<< metal4 >>
rect 2017 -15322 19046 -15257
rect 2017 -15324 4280 -15322
rect 2017 -15560 2354 -15324
rect 2590 -15560 2674 -15324
rect 2910 -15560 2994 -15324
rect 3230 -15558 4280 -15324
rect 4516 -15558 4600 -15322
rect 4836 -15558 4920 -15322
rect 5156 -15324 7668 -15322
rect 5156 -15558 5738 -15324
rect 3230 -15560 5738 -15558
rect 5974 -15560 6058 -15324
rect 6294 -15560 6378 -15324
rect 6614 -15558 7668 -15324
rect 7904 -15558 7988 -15322
rect 8224 -15558 8308 -15322
rect 8544 -15324 11053 -15322
rect 8544 -15558 9123 -15324
rect 6614 -15560 9123 -15558
rect 9359 -15560 9443 -15324
rect 9679 -15560 9763 -15324
rect 9999 -15558 11053 -15324
rect 11289 -15558 11373 -15322
rect 11609 -15558 11693 -15322
rect 11929 -15324 14439 -15322
rect 11929 -15558 12511 -15324
rect 9999 -15560 12511 -15558
rect 12747 -15560 12831 -15324
rect 13067 -15560 13151 -15324
rect 13387 -15558 14439 -15324
rect 14675 -15558 14759 -15322
rect 14995 -15558 15079 -15322
rect 15315 -15324 17825 -15322
rect 15315 -15558 15895 -15324
rect 13387 -15560 15895 -15558
rect 16131 -15560 16215 -15324
rect 16451 -15560 16535 -15324
rect 16771 -15558 17825 -15324
rect 18061 -15558 18145 -15322
rect 18381 -15558 18465 -15322
rect 18701 -15558 19046 -15322
rect 16771 -15560 19046 -15558
rect 2017 -15623 19046 -15560
rect 2194 -17007 5322 -16918
rect 5580 -17007 8708 -16918
rect 8966 -17007 12094 -16918
rect 12352 -17007 15480 -16918
rect 15738 -17007 18866 -16918
rect 2194 -18296 5322 -18207
rect 5580 -18296 8708 -18207
rect 8966 -18296 12094 -18207
rect 12352 -18296 15480 -18207
rect 15738 -18296 18866 -18207
rect 2194 -19585 5322 -19496
rect 5580 -19585 8708 -19496
rect 8966 -19585 12094 -19496
rect 12352 -19585 15480 -19496
rect 15738 -19585 18866 -19496
rect 2194 -20874 5322 -20785
rect 5580 -20874 8708 -20785
rect 8966 -20874 12094 -20785
rect 12352 -20874 15480 -20785
rect 15738 -20874 18866 -20785
rect 2194 -22163 5322 -22074
rect 5580 -22163 8708 -22074
rect 8966 -22163 12094 -22074
rect 12352 -22163 15480 -22074
rect 15738 -22163 18866 -22074
rect 2194 -23452 5322 -23363
rect 5580 -23452 8708 -23363
rect 8966 -23452 12094 -23363
rect 12352 -23452 15480 -23363
rect 15738 -23452 18866 -23363
rect 2194 -24741 5322 -24652
rect 5580 -24741 8708 -24652
rect 8966 -24741 12094 -24652
rect 12352 -24741 15480 -24652
rect 15738 -24741 18866 -24652
<< via4 >>
rect 2354 -15560 2590 -15324
rect 2674 -15560 2910 -15324
rect 2994 -15560 3230 -15324
rect 4280 -15558 4516 -15322
rect 4600 -15558 4836 -15322
rect 4920 -15558 5156 -15322
rect 5738 -15560 5974 -15324
rect 6058 -15560 6294 -15324
rect 6378 -15560 6614 -15324
rect 7668 -15558 7904 -15322
rect 7988 -15558 8224 -15322
rect 8308 -15558 8544 -15322
rect 9123 -15560 9359 -15324
rect 9443 -15560 9679 -15324
rect 9763 -15560 9999 -15324
rect 11053 -15558 11289 -15322
rect 11373 -15558 11609 -15322
rect 11693 -15558 11929 -15322
rect 12511 -15560 12747 -15324
rect 12831 -15560 13067 -15324
rect 13151 -15560 13387 -15324
rect 14439 -15558 14675 -15322
rect 14759 -15558 14995 -15322
rect 15079 -15558 15315 -15322
rect 15895 -15560 16131 -15324
rect 16215 -15560 16451 -15324
rect 16535 -15560 16771 -15324
rect 17825 -15558 18061 -15322
rect 18145 -15558 18381 -15322
rect 18465 -15558 18701 -15322
<< metal5 >>
rect 2310 -15324 3278 -15257
rect 2310 -15560 2354 -15324
rect 2590 -15560 2674 -15324
rect 2910 -15560 2994 -15324
rect 3230 -15560 3278 -15324
rect 2310 -15834 3278 -15560
rect 4238 -15322 5206 -15257
rect 4238 -15558 4280 -15322
rect 4516 -15558 4600 -15322
rect 4836 -15558 4920 -15322
rect 5156 -15558 5206 -15322
rect 4238 -15834 5206 -15558
rect 5696 -15324 6664 -15257
rect 5696 -15560 5738 -15324
rect 5974 -15560 6058 -15324
rect 6294 -15560 6378 -15324
rect 6614 -15560 6664 -15324
rect 5696 -15834 6664 -15560
rect 7624 -15322 8592 -15257
rect 7624 -15558 7668 -15322
rect 7904 -15558 7988 -15322
rect 8224 -15558 8308 -15322
rect 8544 -15558 8592 -15322
rect 7624 -15834 8592 -15558
rect 9082 -15324 10050 -15257
rect 9082 -15560 9123 -15324
rect 9359 -15560 9443 -15324
rect 9679 -15560 9763 -15324
rect 9999 -15560 10050 -15324
rect 9082 -15834 10050 -15560
rect 11010 -15322 11978 -15257
rect 11010 -15558 11053 -15322
rect 11289 -15558 11373 -15322
rect 11609 -15558 11693 -15322
rect 11929 -15558 11978 -15322
rect 11010 -15834 11978 -15558
rect 12468 -15324 13436 -15257
rect 12468 -15560 12511 -15324
rect 12747 -15560 12831 -15324
rect 13067 -15560 13151 -15324
rect 13387 -15560 13436 -15324
rect 12468 -15834 13436 -15560
rect 14396 -15322 15364 -15257
rect 14396 -15558 14439 -15322
rect 14675 -15558 14759 -15322
rect 14995 -15558 15079 -15322
rect 15315 -15558 15364 -15322
rect 14396 -15834 15364 -15558
rect 15854 -15324 16822 -15257
rect 15854 -15560 15895 -15324
rect 16131 -15560 16215 -15324
rect 16451 -15560 16535 -15324
rect 16771 -15560 16822 -15324
rect 15854 -15834 16822 -15560
rect 17782 -15322 18750 -15257
rect 17782 -15558 17825 -15322
rect 18061 -15558 18145 -15322
rect 18381 -15558 18465 -15322
rect 18701 -15558 18750 -15322
rect 17782 -15834 18750 -15558
rect 2310 -17123 3278 -16802
rect 4238 -17123 5206 -16802
rect 5696 -17123 6664 -16802
rect 7624 -17123 8592 -16802
rect 9082 -17123 10050 -16802
rect 11010 -17123 11978 -16802
rect 12468 -17123 13436 -16802
rect 14396 -17123 15364 -16802
rect 15854 -17123 16822 -16802
rect 17782 -17123 18750 -16802
rect 2310 -18412 3278 -18091
rect 4238 -18412 5206 -18091
rect 5696 -18412 6664 -18091
rect 7624 -18412 8592 -18091
rect 9082 -18412 10050 -18091
rect 11010 -18412 11978 -18091
rect 12468 -18412 13436 -18091
rect 14396 -18412 15364 -18091
rect 15854 -18412 16822 -18091
rect 17782 -18412 18750 -18091
rect 2310 -19701 3278 -19380
rect 4238 -19701 5206 -19380
rect 5696 -19701 6664 -19380
rect 7624 -19701 8592 -19380
rect 9082 -19701 10050 -19380
rect 11010 -19701 11978 -19380
rect 12468 -19701 13436 -19380
rect 14396 -19701 15364 -19380
rect 15854 -19701 16822 -19380
rect 17782 -19701 18750 -19380
rect 2310 -20990 3278 -20669
rect 4238 -20990 5206 -20669
rect 5696 -20990 6664 -20669
rect 7624 -20990 8592 -20669
rect 9082 -20990 10050 -20669
rect 11010 -20990 11978 -20669
rect 12468 -20990 13436 -20669
rect 14396 -20990 15364 -20669
rect 15854 -20990 16822 -20669
rect 17782 -20990 18750 -20669
rect 2310 -22279 3278 -21958
rect 4238 -22279 5206 -21958
rect 5696 -22279 6664 -21958
rect 7624 -22279 8592 -21958
rect 9082 -22279 10050 -21958
rect 11010 -22279 11978 -21958
rect 12468 -22279 13436 -21958
rect 14396 -22279 15364 -21958
rect 15854 -22279 16822 -21958
rect 17782 -22279 18750 -21958
rect 2310 -23568 3278 -23247
rect 4238 -23568 5206 -23247
rect 5696 -23568 6664 -23247
rect 7624 -23568 8592 -23247
rect 9082 -23568 10050 -23247
rect 11010 -23568 11978 -23247
rect 12468 -23568 13436 -23247
rect 14396 -23568 15364 -23247
rect 15854 -23568 16822 -23247
rect 17782 -23568 18750 -23247
rect 2310 -24857 3278 -24536
rect 4238 -24857 5206 -24536
rect 5696 -24857 6664 -24536
rect 7624 -24857 8592 -24536
rect 9082 -24857 10050 -24536
rect 11010 -24857 11978 -24536
rect 12468 -24857 13436 -24536
rect 14396 -24857 15364 -24536
rect 15854 -24857 16822 -24536
rect 17782 -24857 18750 -24536
rect 3598 -26158 3918 -25920
rect 6984 -26158 7304 -25920
rect 10370 -26158 10690 -25920
rect 13756 -26158 14076 -25920
rect 17142 -26158 17462 -25920
rect 1997 -26553 19031 -26158
use sky130_fd_pr__cap_mim_m3_1_VCAG9S  sky130_fd_pr__cap_mim_m3_1_VCAG9S_0
array 0 0 1381 0 7 1289
timestamp 1699926577
transform 1 0 18316 0 1 -25341
box -650 -600 731 701
use sky130_fd_pr__cap_mim_m3_1_VCAG9S  sky130_fd_pr__cap_mim_m3_1_VCAG9S_1
array 0 0 -1381 0 7 1289
timestamp 1699926577
transform -1 0 16288 0 1 -25341
box -650 -600 731 701
use sky130_fd_pr__cap_mim_m3_1_VCAG9S  sky130_fd_pr__cap_mim_m3_1_VCAG9S_2
array 0 0 1381 0 7 1289
timestamp 1699926577
transform 1 0 14930 0 1 -25341
box -650 -600 731 701
use sky130_fd_pr__cap_mim_m3_1_VCAG9S  sky130_fd_pr__cap_mim_m3_1_VCAG9S_3
array 0 0 -1381 0 7 1289
timestamp 1699926577
transform -1 0 12902 0 1 -25341
box -650 -600 731 701
use sky130_fd_pr__cap_mim_m3_1_VCAG9S  sky130_fd_pr__cap_mim_m3_1_VCAG9S_4
array 0 0 1381 0 7 1289
timestamp 1699926577
transform 1 0 11544 0 1 -25341
box -650 -600 731 701
use sky130_fd_pr__cap_mim_m3_1_VCAG9S  sky130_fd_pr__cap_mim_m3_1_VCAG9S_5
array 0 0 -1381 0 7 1289
timestamp 1699926577
transform -1 0 9516 0 1 -25341
box -650 -600 731 701
use sky130_fd_pr__cap_mim_m3_1_VCAG9S  sky130_fd_pr__cap_mim_m3_1_VCAG9S_6
array 0 0 1381 0 7 1289
timestamp 1699926577
transform 1 0 8158 0 1 -25341
box -650 -600 731 701
use sky130_fd_pr__cap_mim_m3_1_VCAG9S  sky130_fd_pr__cap_mim_m3_1_VCAG9S_7
array 0 0 -1381 0 7 1289
timestamp 1699926577
transform -1 0 6130 0 1 -25341
box -650 -600 731 701
use sky130_fd_pr__cap_mim_m3_1_VCAG9S  sky130_fd_pr__cap_mim_m3_1_VCAG9S_8
array 0 0 1381 0 7 1289
timestamp 1699926577
transform 1 0 4772 0 1 -25341
box -650 -600 731 701
use sky130_fd_pr__cap_mim_m3_1_VCAG9S  sky130_fd_pr__cap_mim_m3_1_VCAG9S_9
array 0 0 -1381 0 7 1289
timestamp 1699926577
transform -1 0 2744 0 1 -25341
box -650 -600 731 701
use sky130_fd_pr__cap_mim_m3_2_VCAE9S  sky130_fd_pr__cap_mim_m3_2_VCAE9S_0
array 0 0 -1724 0 7 1289
timestamp 1699926577
transform -1 0 18015 0 1 -25341
box -851 -601 873 688
use sky130_fd_pr__cap_mim_m3_2_VCAE9S  sky130_fd_pr__cap_mim_m3_2_VCAE9S_1
array 0 0 1724 0 7 1289
timestamp 1699926577
transform 1 0 16589 0 1 -25341
box -851 -601 873 688
use sky130_fd_pr__cap_mim_m3_2_VCAE9S  sky130_fd_pr__cap_mim_m3_2_VCAE9S_2
array 0 0 -1724 0 7 1289
timestamp 1699926577
transform -1 0 14629 0 1 -25341
box -851 -601 873 688
use sky130_fd_pr__cap_mim_m3_2_VCAE9S  sky130_fd_pr__cap_mim_m3_2_VCAE9S_3
array 0 0 1724 0 7 1289
timestamp 1699926577
transform 1 0 13203 0 1 -25341
box -851 -601 873 688
use sky130_fd_pr__cap_mim_m3_2_VCAE9S  sky130_fd_pr__cap_mim_m3_2_VCAE9S_4
array 0 0 -1724 0 7 1289
timestamp 1699926577
transform -1 0 11243 0 1 -25341
box -851 -601 873 688
use sky130_fd_pr__cap_mim_m3_2_VCAE9S  sky130_fd_pr__cap_mim_m3_2_VCAE9S_5
array 0 0 1724 0 7 1289
timestamp 1699926577
transform 1 0 9817 0 1 -25341
box -851 -601 873 688
use sky130_fd_pr__cap_mim_m3_2_VCAE9S  sky130_fd_pr__cap_mim_m3_2_VCAE9S_6
array 0 0 -1724 0 7 1289
timestamp 1699926577
transform -1 0 7857 0 1 -25341
box -851 -601 873 688
use sky130_fd_pr__cap_mim_m3_2_VCAE9S  sky130_fd_pr__cap_mim_m3_2_VCAE9S_7
array 0 0 1724 0 7 1289
timestamp 1699926577
transform 1 0 6431 0 1 -25341
box -851 -601 873 688
use sky130_fd_pr__cap_mim_m3_2_VCAE9S  sky130_fd_pr__cap_mim_m3_2_VCAE9S_8
array 0 0 -1724 0 7 1289
timestamp 1699926577
transform -1 0 4471 0 1 -25341
box -851 -601 873 688
use sky130_fd_pr__cap_mim_m3_2_VCAE9S  XC2
array 0 0 1724 0 7 1289
timestamp 1699926577
transform 1 0 3045 0 1 -25341
box -851 -601 873 688
<< labels >>
flabel metal4 s 3664 -15423 3664 -15423 0 FreeSans 25 0 0 0 vss
flabel metal5 s 3731 -26364 3731 -26364 0 FreeSans 25 0 0 0 holdval
<< end >>
