magic
tech sky130A
magscale 1 2
timestamp 1693827120
<< metal2 >>
rect -2079 78 1 100
rect -2079 22 -2044 78
rect -1988 22 -1964 78
rect -1908 22 -1884 78
rect -1828 22 -1804 78
rect -1748 22 -1724 78
rect -1668 22 -1644 78
rect -1588 22 -1564 78
rect -1508 22 -1484 78
rect -1428 22 -1404 78
rect -1348 22 -1324 78
rect -1268 22 -1244 78
rect -1188 22 -1164 78
rect -1108 22 -1084 78
rect -1028 22 -1004 78
rect -948 22 -924 78
rect -868 22 -844 78
rect -788 22 -764 78
rect -708 22 -684 78
rect -628 22 -604 78
rect -548 22 -524 78
rect -468 22 -444 78
rect -388 22 -364 78
rect -308 22 -284 78
rect -228 22 -204 78
rect -148 22 -124 78
rect -68 22 1 78
rect -2079 0 1 22
<< via2 >>
rect -2044 22 -1988 78
rect -1964 22 -1908 78
rect -1884 22 -1828 78
rect -1804 22 -1748 78
rect -1724 22 -1668 78
rect -1644 22 -1588 78
rect -1564 22 -1508 78
rect -1484 22 -1428 78
rect -1404 22 -1348 78
rect -1324 22 -1268 78
rect -1244 22 -1188 78
rect -1164 22 -1108 78
rect -1084 22 -1028 78
rect -1004 22 -948 78
rect -924 22 -868 78
rect -844 22 -788 78
rect -764 22 -708 78
rect -684 22 -628 78
rect -604 22 -548 78
rect -524 22 -468 78
rect -444 22 -388 78
rect -364 22 -308 78
rect -284 22 -228 78
rect -204 22 -148 78
rect -124 22 -68 78
<< metal3 >>
rect -2079 78 1 100
rect -2079 22 -2044 78
rect -1988 22 -1964 78
rect -1908 22 -1884 78
rect -1828 22 -1804 78
rect -1748 22 -1724 78
rect -1668 22 -1644 78
rect -1588 22 -1564 78
rect -1508 22 -1484 78
rect -1428 22 -1404 78
rect -1348 22 -1324 78
rect -1268 22 -1244 78
rect -1188 22 -1164 78
rect -1108 22 -1084 78
rect -1028 22 -1004 78
rect -948 22 -924 78
rect -868 22 -844 78
rect -788 22 -764 78
rect -708 22 -684 78
rect -628 22 -604 78
rect -548 22 -524 78
rect -468 22 -444 78
rect -388 22 -364 78
rect -308 22 -284 78
rect -228 22 -204 78
rect -148 22 -124 78
rect -68 22 1 78
rect -2079 0 1 22
<< end >>
