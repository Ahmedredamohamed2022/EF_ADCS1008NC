magic
tech sky130A
magscale 1 2
timestamp 1693827120
<< metal3 >>
rect -1186 992 1186 1040
rect -1186 928 1102 992
rect 1166 928 1186 992
rect -1186 912 1186 928
rect -1186 848 1102 912
rect 1166 848 1186 912
rect -1186 832 1186 848
rect -1186 768 1102 832
rect 1166 768 1186 832
rect -1186 752 1186 768
rect -1186 688 1102 752
rect 1166 688 1186 752
rect -1186 672 1186 688
rect -1186 608 1102 672
rect 1166 608 1186 672
rect -1186 592 1186 608
rect -1186 528 1102 592
rect 1166 528 1186 592
rect -1186 512 1186 528
rect -1186 448 1102 512
rect 1166 448 1186 512
rect -1186 432 1186 448
rect -1186 368 1102 432
rect 1166 368 1186 432
rect -1186 352 1186 368
rect -1186 288 1102 352
rect 1166 288 1186 352
rect -1186 272 1186 288
rect -1186 208 1102 272
rect 1166 208 1186 272
rect -1186 192 1186 208
rect -1186 128 1102 192
rect 1166 128 1186 192
rect -1186 112 1186 128
rect -1186 48 1102 112
rect 1166 48 1186 112
rect -1186 32 1186 48
rect -1186 -32 1102 32
rect 1166 -32 1186 32
rect -1186 -48 1186 -32
rect -1186 -112 1102 -48
rect 1166 -112 1186 -48
rect -1186 -128 1186 -112
rect -1186 -192 1102 -128
rect 1166 -192 1186 -128
rect -1186 -208 1186 -192
rect -1186 -272 1102 -208
rect 1166 -272 1186 -208
rect -1186 -288 1186 -272
rect -1186 -352 1102 -288
rect 1166 -352 1186 -288
rect -1186 -368 1186 -352
rect -1186 -432 1102 -368
rect 1166 -432 1186 -368
rect -1186 -448 1186 -432
rect -1186 -512 1102 -448
rect 1166 -512 1186 -448
rect -1186 -528 1186 -512
rect -1186 -592 1102 -528
rect 1166 -592 1186 -528
rect -1186 -608 1186 -592
rect -1186 -672 1102 -608
rect 1166 -672 1186 -608
rect -1186 -688 1186 -672
rect -1186 -752 1102 -688
rect 1166 -752 1186 -688
rect -1186 -768 1186 -752
rect -1186 -832 1102 -768
rect 1166 -832 1186 -768
rect -1186 -848 1186 -832
rect -1186 -912 1102 -848
rect 1166 -912 1186 -848
rect -1186 -928 1186 -912
rect -1186 -992 1102 -928
rect 1166 -992 1186 -928
rect -1186 -1040 1186 -992
<< via3 >>
rect 1102 928 1166 992
rect 1102 848 1166 912
rect 1102 768 1166 832
rect 1102 688 1166 752
rect 1102 608 1166 672
rect 1102 528 1166 592
rect 1102 448 1166 512
rect 1102 368 1166 432
rect 1102 288 1166 352
rect 1102 208 1166 272
rect 1102 128 1166 192
rect 1102 48 1166 112
rect 1102 -32 1166 32
rect 1102 -112 1166 -48
rect 1102 -192 1166 -128
rect 1102 -272 1166 -208
rect 1102 -352 1166 -288
rect 1102 -432 1166 -368
rect 1102 -512 1166 -448
rect 1102 -592 1166 -528
rect 1102 -672 1166 -608
rect 1102 -752 1166 -688
rect 1102 -832 1166 -768
rect 1102 -912 1166 -848
rect 1102 -992 1166 -928
<< mimcap >>
rect -1146 952 854 1000
rect -1146 -952 -1098 952
rect 806 -952 854 952
rect -1146 -1000 854 -952
<< mimcapcontact >>
rect -1098 -952 806 952
<< metal4 >>
rect 1086 992 1182 1028
rect -1107 952 815 961
rect -1107 -952 -1098 952
rect 806 -952 815 952
rect -1107 -961 815 -952
rect 1086 928 1102 992
rect 1166 928 1182 992
rect 1086 912 1182 928
rect 1086 848 1102 912
rect 1166 848 1182 912
rect 1086 832 1182 848
rect 1086 768 1102 832
rect 1166 768 1182 832
rect 1086 752 1182 768
rect 1086 688 1102 752
rect 1166 688 1182 752
rect 1086 672 1182 688
rect 1086 608 1102 672
rect 1166 608 1182 672
rect 1086 592 1182 608
rect 1086 528 1102 592
rect 1166 528 1182 592
rect 1086 512 1182 528
rect 1086 448 1102 512
rect 1166 448 1182 512
rect 1086 432 1182 448
rect 1086 368 1102 432
rect 1166 368 1182 432
rect 1086 352 1182 368
rect 1086 288 1102 352
rect 1166 288 1182 352
rect 1086 272 1182 288
rect 1086 208 1102 272
rect 1166 208 1182 272
rect 1086 192 1182 208
rect 1086 128 1102 192
rect 1166 128 1182 192
rect 1086 112 1182 128
rect 1086 48 1102 112
rect 1166 48 1182 112
rect 1086 32 1182 48
rect 1086 -32 1102 32
rect 1166 -32 1182 32
rect 1086 -48 1182 -32
rect 1086 -112 1102 -48
rect 1166 -112 1182 -48
rect 1086 -128 1182 -112
rect 1086 -192 1102 -128
rect 1166 -192 1182 -128
rect 1086 -208 1182 -192
rect 1086 -272 1102 -208
rect 1166 -272 1182 -208
rect 1086 -288 1182 -272
rect 1086 -352 1102 -288
rect 1166 -352 1182 -288
rect 1086 -368 1182 -352
rect 1086 -432 1102 -368
rect 1166 -432 1182 -368
rect 1086 -448 1182 -432
rect 1086 -512 1102 -448
rect 1166 -512 1182 -448
rect 1086 -528 1182 -512
rect 1086 -592 1102 -528
rect 1166 -592 1182 -528
rect 1086 -608 1182 -592
rect 1086 -672 1102 -608
rect 1166 -672 1182 -608
rect 1086 -688 1182 -672
rect 1086 -752 1102 -688
rect 1166 -752 1182 -688
rect 1086 -768 1182 -752
rect 1086 -832 1102 -768
rect 1166 -832 1182 -768
rect 1086 -848 1182 -832
rect 1086 -912 1102 -848
rect 1166 -912 1182 -848
rect 1086 -928 1182 -912
rect 1086 -992 1102 -928
rect 1166 -992 1182 -928
rect 1086 -1028 1182 -992
<< properties >>
string FIXED_BBOX -1186 -1040 894 1040
<< end >>
