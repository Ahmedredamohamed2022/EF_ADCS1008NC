magic
tech sky130A
magscale 1 2
timestamp 1699926577
<< metal3 >>
rect -2486 2312 2486 2340
rect -2486 2248 2402 2312
rect 2466 2248 2486 2312
rect -2486 2232 2486 2248
rect -2486 2168 2402 2232
rect 2466 2168 2486 2232
rect -2486 2152 2486 2168
rect -2486 2088 2402 2152
rect 2466 2088 2486 2152
rect -2486 2072 2486 2088
rect -2486 2008 2402 2072
rect 2466 2008 2486 2072
rect -2486 1992 2486 2008
rect -2486 1928 2402 1992
rect 2466 1928 2486 1992
rect -2486 1912 2486 1928
rect -2486 1848 2402 1912
rect 2466 1848 2486 1912
rect -2486 1832 2486 1848
rect -2486 1768 2402 1832
rect 2466 1768 2486 1832
rect -2486 1752 2486 1768
rect -2486 1688 2402 1752
rect 2466 1688 2486 1752
rect -2486 1672 2486 1688
rect -2486 1608 2402 1672
rect 2466 1608 2486 1672
rect -2486 1592 2486 1608
rect -2486 1528 2402 1592
rect 2466 1528 2486 1592
rect -2486 1512 2486 1528
rect -2486 1448 2402 1512
rect 2466 1448 2486 1512
rect -2486 1432 2486 1448
rect -2486 1368 2402 1432
rect 2466 1368 2486 1432
rect -2486 1352 2486 1368
rect -2486 1288 2402 1352
rect 2466 1288 2486 1352
rect -2486 1272 2486 1288
rect -2486 1208 2402 1272
rect 2466 1208 2486 1272
rect -2486 1192 2486 1208
rect -2486 1128 2402 1192
rect 2466 1128 2486 1192
rect -2486 1112 2486 1128
rect -2486 1048 2402 1112
rect 2466 1048 2486 1112
rect -2486 1032 2486 1048
rect -2486 968 2402 1032
rect 2466 968 2486 1032
rect -2486 952 2486 968
rect -2486 888 2402 952
rect 2466 888 2486 952
rect -2486 872 2486 888
rect -2486 808 2402 872
rect 2466 808 2486 872
rect -2486 792 2486 808
rect -2486 728 2402 792
rect 2466 728 2486 792
rect -2486 712 2486 728
rect -2486 648 2402 712
rect 2466 648 2486 712
rect -2486 632 2486 648
rect -2486 568 2402 632
rect 2466 568 2486 632
rect -2486 552 2486 568
rect -2486 488 2402 552
rect 2466 488 2486 552
rect -2486 472 2486 488
rect -2486 408 2402 472
rect 2466 408 2486 472
rect -2486 392 2486 408
rect -2486 328 2402 392
rect 2466 328 2486 392
rect -2486 312 2486 328
rect -2486 248 2402 312
rect 2466 248 2486 312
rect -2486 232 2486 248
rect -2486 168 2402 232
rect 2466 168 2486 232
rect -2486 152 2486 168
rect -2486 88 2402 152
rect 2466 88 2486 152
rect -2486 72 2486 88
rect -2486 8 2402 72
rect 2466 8 2486 72
rect -2486 -8 2486 8
rect -2486 -72 2402 -8
rect 2466 -72 2486 -8
rect -2486 -88 2486 -72
rect -2486 -152 2402 -88
rect 2466 -152 2486 -88
rect -2486 -168 2486 -152
rect -2486 -232 2402 -168
rect 2466 -232 2486 -168
rect -2486 -248 2486 -232
rect -2486 -312 2402 -248
rect 2466 -312 2486 -248
rect -2486 -328 2486 -312
rect -2486 -392 2402 -328
rect 2466 -392 2486 -328
rect -2486 -408 2486 -392
rect -2486 -472 2402 -408
rect 2466 -472 2486 -408
rect -2486 -488 2486 -472
rect -2486 -552 2402 -488
rect 2466 -552 2486 -488
rect -2486 -568 2486 -552
rect -2486 -632 2402 -568
rect 2466 -632 2486 -568
rect -2486 -648 2486 -632
rect -2486 -712 2402 -648
rect 2466 -712 2486 -648
rect -2486 -728 2486 -712
rect -2486 -792 2402 -728
rect 2466 -792 2486 -728
rect -2486 -808 2486 -792
rect -2486 -872 2402 -808
rect 2466 -872 2486 -808
rect -2486 -888 2486 -872
rect -2486 -952 2402 -888
rect 2466 -952 2486 -888
rect -2486 -968 2486 -952
rect -2486 -1032 2402 -968
rect 2466 -1032 2486 -968
rect -2486 -1048 2486 -1032
rect -2486 -1112 2402 -1048
rect 2466 -1112 2486 -1048
rect -2486 -1128 2486 -1112
rect -2486 -1192 2402 -1128
rect 2466 -1192 2486 -1128
rect -2486 -1208 2486 -1192
rect -2486 -1272 2402 -1208
rect 2466 -1272 2486 -1208
rect -2486 -1288 2486 -1272
rect -2486 -1352 2402 -1288
rect 2466 -1352 2486 -1288
rect -2486 -1368 2486 -1352
rect -2486 -1432 2402 -1368
rect 2466 -1432 2486 -1368
rect -2486 -1448 2486 -1432
rect -2486 -1512 2402 -1448
rect 2466 -1512 2486 -1448
rect -2486 -1528 2486 -1512
rect -2486 -1592 2402 -1528
rect 2466 -1592 2486 -1528
rect -2486 -1608 2486 -1592
rect -2486 -1672 2402 -1608
rect 2466 -1672 2486 -1608
rect -2486 -1688 2486 -1672
rect -2486 -1752 2402 -1688
rect 2466 -1752 2486 -1688
rect -2486 -1768 2486 -1752
rect -2486 -1832 2402 -1768
rect 2466 -1832 2486 -1768
rect -2486 -1848 2486 -1832
rect -2486 -1912 2402 -1848
rect 2466 -1912 2486 -1848
rect -2486 -1928 2486 -1912
rect -2486 -1992 2402 -1928
rect 2466 -1992 2486 -1928
rect -2486 -2008 2486 -1992
rect -2486 -2072 2402 -2008
rect 2466 -2072 2486 -2008
rect -2486 -2088 2486 -2072
rect -2486 -2152 2402 -2088
rect 2466 -2152 2486 -2088
rect -2486 -2168 2486 -2152
rect -2486 -2232 2402 -2168
rect 2466 -2232 2486 -2168
rect -2486 -2248 2486 -2232
rect -2486 -2312 2402 -2248
rect 2466 -2312 2486 -2248
rect -2486 -2340 2486 -2312
<< via3 >>
rect 2402 2248 2466 2312
rect 2402 2168 2466 2232
rect 2402 2088 2466 2152
rect 2402 2008 2466 2072
rect 2402 1928 2466 1992
rect 2402 1848 2466 1912
rect 2402 1768 2466 1832
rect 2402 1688 2466 1752
rect 2402 1608 2466 1672
rect 2402 1528 2466 1592
rect 2402 1448 2466 1512
rect 2402 1368 2466 1432
rect 2402 1288 2466 1352
rect 2402 1208 2466 1272
rect 2402 1128 2466 1192
rect 2402 1048 2466 1112
rect 2402 968 2466 1032
rect 2402 888 2466 952
rect 2402 808 2466 872
rect 2402 728 2466 792
rect 2402 648 2466 712
rect 2402 568 2466 632
rect 2402 488 2466 552
rect 2402 408 2466 472
rect 2402 328 2466 392
rect 2402 248 2466 312
rect 2402 168 2466 232
rect 2402 88 2466 152
rect 2402 8 2466 72
rect 2402 -72 2466 -8
rect 2402 -152 2466 -88
rect 2402 -232 2466 -168
rect 2402 -312 2466 -248
rect 2402 -392 2466 -328
rect 2402 -472 2466 -408
rect 2402 -552 2466 -488
rect 2402 -632 2466 -568
rect 2402 -712 2466 -648
rect 2402 -792 2466 -728
rect 2402 -872 2466 -808
rect 2402 -952 2466 -888
rect 2402 -1032 2466 -968
rect 2402 -1112 2466 -1048
rect 2402 -1192 2466 -1128
rect 2402 -1272 2466 -1208
rect 2402 -1352 2466 -1288
rect 2402 -1432 2466 -1368
rect 2402 -1512 2466 -1448
rect 2402 -1592 2466 -1528
rect 2402 -1672 2466 -1608
rect 2402 -1752 2466 -1688
rect 2402 -1832 2466 -1768
rect 2402 -1912 2466 -1848
rect 2402 -1992 2466 -1928
rect 2402 -2072 2466 -2008
rect 2402 -2152 2466 -2088
rect 2402 -2232 2466 -2168
rect 2402 -2312 2466 -2248
<< mimcap >>
rect -2446 2232 2154 2300
rect -2446 -2232 -2378 2232
rect 2086 -2232 2154 2232
rect -2446 -2300 2154 -2232
<< mimcapcontact >>
rect -2378 -2232 2086 2232
<< metal4 >>
rect 2386 2312 2482 2328
rect -2407 2232 2115 2261
rect -2407 -2232 -2378 2232
rect 2086 -2232 2115 2232
rect -2407 -2261 2115 -2232
rect 2386 2248 2402 2312
rect 2466 2248 2482 2312
rect 2386 2232 2482 2248
rect 2386 2168 2402 2232
rect 2466 2168 2482 2232
rect 2386 2152 2482 2168
rect 2386 2088 2402 2152
rect 2466 2088 2482 2152
rect 2386 2072 2482 2088
rect 2386 2008 2402 2072
rect 2466 2008 2482 2072
rect 2386 1992 2482 2008
rect 2386 1928 2402 1992
rect 2466 1928 2482 1992
rect 2386 1912 2482 1928
rect 2386 1848 2402 1912
rect 2466 1848 2482 1912
rect 2386 1832 2482 1848
rect 2386 1768 2402 1832
rect 2466 1768 2482 1832
rect 2386 1752 2482 1768
rect 2386 1688 2402 1752
rect 2466 1688 2482 1752
rect 2386 1672 2482 1688
rect 2386 1608 2402 1672
rect 2466 1608 2482 1672
rect 2386 1592 2482 1608
rect 2386 1528 2402 1592
rect 2466 1528 2482 1592
rect 2386 1512 2482 1528
rect 2386 1448 2402 1512
rect 2466 1448 2482 1512
rect 2386 1432 2482 1448
rect 2386 1368 2402 1432
rect 2466 1368 2482 1432
rect 2386 1352 2482 1368
rect 2386 1288 2402 1352
rect 2466 1288 2482 1352
rect 2386 1272 2482 1288
rect 2386 1208 2402 1272
rect 2466 1208 2482 1272
rect 2386 1192 2482 1208
rect 2386 1128 2402 1192
rect 2466 1128 2482 1192
rect 2386 1112 2482 1128
rect 2386 1048 2402 1112
rect 2466 1048 2482 1112
rect 2386 1032 2482 1048
rect 2386 968 2402 1032
rect 2466 968 2482 1032
rect 2386 952 2482 968
rect 2386 888 2402 952
rect 2466 888 2482 952
rect 2386 872 2482 888
rect 2386 808 2402 872
rect 2466 808 2482 872
rect 2386 792 2482 808
rect 2386 728 2402 792
rect 2466 728 2482 792
rect 2386 712 2482 728
rect 2386 648 2402 712
rect 2466 648 2482 712
rect 2386 632 2482 648
rect 2386 568 2402 632
rect 2466 568 2482 632
rect 2386 552 2482 568
rect 2386 488 2402 552
rect 2466 488 2482 552
rect 2386 472 2482 488
rect 2386 408 2402 472
rect 2466 408 2482 472
rect 2386 392 2482 408
rect 2386 328 2402 392
rect 2466 328 2482 392
rect 2386 312 2482 328
rect 2386 248 2402 312
rect 2466 248 2482 312
rect 2386 232 2482 248
rect 2386 168 2402 232
rect 2466 168 2482 232
rect 2386 152 2482 168
rect 2386 88 2402 152
rect 2466 88 2482 152
rect 2386 72 2482 88
rect 2386 8 2402 72
rect 2466 8 2482 72
rect 2386 -8 2482 8
rect 2386 -72 2402 -8
rect 2466 -72 2482 -8
rect 2386 -88 2482 -72
rect 2386 -152 2402 -88
rect 2466 -152 2482 -88
rect 2386 -168 2482 -152
rect 2386 -232 2402 -168
rect 2466 -232 2482 -168
rect 2386 -248 2482 -232
rect 2386 -312 2402 -248
rect 2466 -312 2482 -248
rect 2386 -328 2482 -312
rect 2386 -392 2402 -328
rect 2466 -392 2482 -328
rect 2386 -408 2482 -392
rect 2386 -472 2402 -408
rect 2466 -472 2482 -408
rect 2386 -488 2482 -472
rect 2386 -552 2402 -488
rect 2466 -552 2482 -488
rect 2386 -568 2482 -552
rect 2386 -632 2402 -568
rect 2466 -632 2482 -568
rect 2386 -648 2482 -632
rect 2386 -712 2402 -648
rect 2466 -712 2482 -648
rect 2386 -728 2482 -712
rect 2386 -792 2402 -728
rect 2466 -792 2482 -728
rect 2386 -808 2482 -792
rect 2386 -872 2402 -808
rect 2466 -872 2482 -808
rect 2386 -888 2482 -872
rect 2386 -952 2402 -888
rect 2466 -952 2482 -888
rect 2386 -968 2482 -952
rect 2386 -1032 2402 -968
rect 2466 -1032 2482 -968
rect 2386 -1048 2482 -1032
rect 2386 -1112 2402 -1048
rect 2466 -1112 2482 -1048
rect 2386 -1128 2482 -1112
rect 2386 -1192 2402 -1128
rect 2466 -1192 2482 -1128
rect 2386 -1208 2482 -1192
rect 2386 -1272 2402 -1208
rect 2466 -1272 2482 -1208
rect 2386 -1288 2482 -1272
rect 2386 -1352 2402 -1288
rect 2466 -1352 2482 -1288
rect 2386 -1368 2482 -1352
rect 2386 -1432 2402 -1368
rect 2466 -1432 2482 -1368
rect 2386 -1448 2482 -1432
rect 2386 -1512 2402 -1448
rect 2466 -1512 2482 -1448
rect 2386 -1528 2482 -1512
rect 2386 -1592 2402 -1528
rect 2466 -1592 2482 -1528
rect 2386 -1608 2482 -1592
rect 2386 -1672 2402 -1608
rect 2466 -1672 2482 -1608
rect 2386 -1688 2482 -1672
rect 2386 -1752 2402 -1688
rect 2466 -1752 2482 -1688
rect 2386 -1768 2482 -1752
rect 2386 -1832 2402 -1768
rect 2466 -1832 2482 -1768
rect 2386 -1848 2482 -1832
rect 2386 -1912 2402 -1848
rect 2466 -1912 2482 -1848
rect 2386 -1928 2482 -1912
rect 2386 -1992 2402 -1928
rect 2466 -1992 2482 -1928
rect 2386 -2008 2482 -1992
rect 2386 -2072 2402 -2008
rect 2466 -2072 2482 -2008
rect 2386 -2088 2482 -2072
rect 2386 -2152 2402 -2088
rect 2466 -2152 2482 -2088
rect 2386 -2168 2482 -2152
rect 2386 -2232 2402 -2168
rect 2466 -2232 2482 -2168
rect 2386 -2248 2482 -2232
rect 2386 -2312 2402 -2248
rect 2466 -2312 2482 -2248
rect 2386 -2328 2482 -2312
<< properties >>
string FIXED_BBOX -2486 -2340 2194 2340
<< end >>
