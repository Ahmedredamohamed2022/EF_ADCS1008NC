VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO EF_ADCS1008NC
  CLASS BLOCK ;
  FOREIGN EF_ADCS1008NC ;
  ORIGIN 7.750 460.805 ;
  SIZE 345.570 BY 525.835 ;
  PIN B[0]
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 168.510 34.080 170.050 34.380 ;
    END
  END B[0]
  PIN B[1]
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 168.500 33.390 170.040 33.690 ;
    END
  END B[1]
  PIN B[2]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 168.520 32.720 170.060 33.020 ;
    END
  END B[2]
  PIN VIN[0]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 133.760 63.490 134.215 64.980 ;
    END
  END VIN[0]
  PIN VIN[1]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 116.540 63.490 117.020 65.000 ;
    END
  END VIN[1]
  PIN VIN[2]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 100.020 63.510 100.500 65.020 ;
    END
  END VIN[2]
  PIN VIN[3]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 83.140 63.530 83.600 65.010 ;
    END
  END VIN[3]
  PIN VIN[4]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 66.590 63.500 67.050 64.980 ;
    END
  END VIN[4]
  PIN VIN[5]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 50.070 63.510 50.530 64.990 ;
    END
  END VIN[5]
  PIN VIN[6]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 33.080 63.510 33.540 64.990 ;
    END
  END VIN[6]
  PIN VIN[7]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 16.090 63.530 16.550 65.010 ;
    END
  END VIN[7]
  PIN HOLD
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.360000 ;
    PORT
      LAYER met3 ;
        RECT -6.040 -18.730 -2.890 -17.720 ;
    END
    PORT
      LAYER met1 ;
        RECT -0.180 -18.745 0.820 -17.745 ;
    END
  END HOLD
  PIN CMP
    ANTENNADIFFAREA 0.492900 ;
    PORT
      LAYER met3 ;
        RECT 167.940 -42.450 170.010 -41.460 ;
    END
  END CMP
  PIN DATA[9]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -0.030 -132.980 5.730 -132.100 ;
    END
  END DATA[9]
  PIN DATA[8]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -0.010 -166.610 5.750 -165.730 ;
    END
  END DATA[8]
  PIN DATA[7]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -0.050 -200.190 5.710 -199.310 ;
    END
  END DATA[7]
  PIN DATA[6]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.010 -233.660 5.770 -232.780 ;
    END
  END DATA[6]
  PIN DATA[5]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.030 -267.510 5.790 -266.630 ;
    END
  END DATA[5]
  PIN DATA[0]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -0.030 -302.440 5.730 -301.560 ;
    END
  END DATA[0]
  PIN DATA[1]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT 0.010 -335.970 5.770 -335.090 ;
    END
  END DATA[1]
  PIN DATA[2]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -0.010 -369.570 5.750 -368.690 ;
    END
  END DATA[2]
  PIN DATA[3]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -0.050 -403.080 5.710 -402.200 ;
    END
  END DATA[3]
  PIN DATA[4]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -0.030 -436.970 5.730 -436.090 ;
    END
  END DATA[4]
  PIN VH
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met3 ;
        RECT -0.030 -272.070 5.730 -271.190 ;
    END
  END VH
  PIN VL
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met3 ;
        RECT -0.080 -274.400 5.680 -273.520 ;
    END
  END VL
  PIN RST
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER met3 ;
        RECT -2.030 -75.430 2.070 -74.420 ;
    END
  END RST
  PIN DVDD
    ANTENNAGATEAREA 47.261497 ;
    ANTENNADIFFAREA 93.596451 ;
    PORT
      LAYER met3 ;
        RECT 0.010 -444.670 7.200 -442.680 ;
    END
  END DVDD
  PIN DVSS
    ANTENNAGATEAREA 74.759102 ;
    ANTENNADIFFAREA 1023.766663 ;
    PORT
      LAYER met3 ;
        RECT -0.020 -447.340 7.170 -445.350 ;
    END
  END DVSS
  PIN VSS
    ANTENNAGATEAREA 130.500000 ;
    ANTENNADIFFAREA 621.362671 ;
    PORT
      LAYER met3 ;
        RECT -0.030 -452.560 7.380 -450.660 ;
    END
  END VSS
  PIN VDD
    ANTENNAGATEAREA 100.000000 ;
    ANTENNADIFFAREA 2509.495605 ;
    PORT
      LAYER met3 ;
        RECT 0.090 -449.800 7.390 -447.860 ;
    END
  END VDD
  PIN EN
    ANTENNAGATEAREA 1.752000 ;
    ANTENNADIFFAREA 1.080000 ;
    PORT
      LAYER met3 ;
        RECT -6.040 -39.960 -3.250 -39.030 ;
    END
  END EN
  OBS
      LAYER li1 ;
        RECT 1.185 -438.520 241.870 54.795 ;
      LAYER met1 ;
        RECT -5.995 -17.465 242.565 55.000 ;
        RECT -5.995 -19.025 -0.460 -17.465 ;
        RECT 1.100 -19.025 242.565 -17.465 ;
        RECT -5.995 -440.835 242.565 -19.025 ;
      LAYER met2 ;
        RECT -6.040 63.250 15.810 65.030 ;
        RECT 16.830 63.250 32.800 65.030 ;
        RECT -6.040 63.230 32.800 63.250 ;
        RECT 33.820 63.230 49.790 65.030 ;
        RECT 50.810 63.230 66.310 65.030 ;
        RECT -6.040 63.220 66.310 63.230 ;
        RECT 67.330 63.250 82.860 65.030 ;
        RECT 83.880 63.250 99.740 65.030 ;
        RECT 67.330 63.230 99.740 63.250 ;
        RECT 100.780 63.230 116.260 65.030 ;
        RECT 67.330 63.220 116.260 63.230 ;
        RECT -6.040 63.210 116.260 63.220 ;
        RECT 117.300 63.210 133.480 65.030 ;
        RECT 134.495 63.210 240.250 65.030 ;
        RECT -6.040 -440.835 240.250 63.210 ;
      LAYER met3 ;
        RECT -6.050 34.780 337.820 63.000 ;
        RECT -6.050 34.090 168.110 34.780 ;
        RECT -6.050 32.990 168.100 34.090 ;
        RECT 170.450 33.680 337.820 34.780 ;
        RECT 170.440 33.420 337.820 33.680 ;
        RECT -6.050 32.320 168.120 32.990 ;
        RECT 170.460 32.320 337.820 33.420 ;
        RECT -6.050 -17.320 337.820 32.320 ;
        RECT -2.490 -19.130 337.820 -17.320 ;
        RECT -6.050 -38.630 337.820 -19.130 ;
        RECT -2.850 -40.360 337.820 -38.630 ;
        RECT -6.050 -41.060 337.820 -40.360 ;
        RECT -6.050 -42.850 167.540 -41.060 ;
        RECT 170.410 -42.850 337.820 -41.060 ;
        RECT -6.050 -74.020 337.820 -42.850 ;
        RECT -6.050 -75.830 -2.430 -74.020 ;
        RECT 2.470 -75.830 337.820 -74.020 ;
        RECT -6.050 -131.700 337.820 -75.830 ;
        RECT -6.050 -133.380 -0.430 -131.700 ;
        RECT 6.130 -133.380 337.820 -131.700 ;
        RECT -6.050 -165.330 337.820 -133.380 ;
        RECT -6.050 -167.010 -0.410 -165.330 ;
        RECT 6.150 -167.010 337.820 -165.330 ;
        RECT -6.050 -198.910 337.820 -167.010 ;
        RECT -6.050 -200.590 -0.450 -198.910 ;
        RECT 6.110 -200.590 337.820 -198.910 ;
        RECT -6.050 -232.380 337.820 -200.590 ;
        RECT -6.050 -234.060 -0.390 -232.380 ;
        RECT 6.170 -234.060 337.820 -232.380 ;
        RECT -6.050 -266.230 337.820 -234.060 ;
        RECT -6.050 -267.910 -0.370 -266.230 ;
        RECT 6.190 -267.910 337.820 -266.230 ;
        RECT -6.050 -270.790 337.820 -267.910 ;
        RECT -6.050 -272.470 -0.430 -270.790 ;
        RECT 6.130 -272.470 337.820 -270.790 ;
        RECT -6.050 -273.120 337.820 -272.470 ;
        RECT -6.050 -274.800 -0.480 -273.120 ;
        RECT 6.080 -274.800 337.820 -273.120 ;
        RECT -6.050 -301.160 337.820 -274.800 ;
        RECT -6.050 -302.840 -0.430 -301.160 ;
        RECT 6.130 -302.840 337.820 -301.160 ;
        RECT -6.050 -334.690 337.820 -302.840 ;
        RECT -6.050 -336.370 -0.390 -334.690 ;
        RECT 6.170 -336.370 337.820 -334.690 ;
        RECT -6.050 -368.290 337.820 -336.370 ;
        RECT -6.050 -369.970 -0.410 -368.290 ;
        RECT 6.150 -369.970 337.820 -368.290 ;
        RECT -6.050 -401.800 337.820 -369.970 ;
        RECT -6.050 -403.480 -0.450 -401.800 ;
        RECT 6.110 -403.480 337.820 -401.800 ;
        RECT -6.050 -435.690 337.820 -403.480 ;
        RECT -6.050 -437.370 -0.430 -435.690 ;
        RECT 6.130 -437.370 337.820 -435.690 ;
        RECT -6.050 -442.280 337.820 -437.370 ;
        RECT -6.050 -444.950 -0.390 -442.280 ;
        RECT -6.050 -447.740 -0.420 -444.950 ;
        RECT 7.600 -445.070 337.820 -442.280 ;
        RECT 7.570 -447.460 337.820 -445.070 ;
        RECT -6.050 -450.200 -0.310 -447.740 ;
        RECT 7.790 -450.200 337.820 -447.460 ;
        RECT -6.050 -450.260 337.820 -450.200 ;
        RECT -6.050 -452.595 -0.430 -450.260 ;
        RECT 7.780 -452.595 337.820 -450.260 ;
      LAYER met4 ;
        RECT -2.170 -452.595 337.650 63.000 ;
      LAYER met5 ;
        RECT 10.895 -68.115 164.925 54.315 ;
  END
END EF_ADCS1008NC
END LIBRARY

