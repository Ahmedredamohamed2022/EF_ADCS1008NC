magic
tech sky130A
magscale 1 2
timestamp 1699926577
<< pwell >>
rect -173 -173 173 173
<< psubdiff >>
rect -147 113 -51 147
rect -17 113 17 147
rect 51 113 147 147
rect -147 51 -113 113
rect 113 51 147 113
rect -147 -17 -113 17
rect 113 -17 147 17
rect -147 -113 -113 -51
rect 113 -113 147 -51
rect -147 -147 -51 -113
rect -17 -147 17 -113
rect 51 -147 147 -113
<< psubdiffcont >>
rect -51 113 -17 147
rect 17 113 51 147
rect -147 17 -113 51
rect -147 -51 -113 -17
rect 113 17 147 51
rect 113 -51 147 -17
rect -51 -147 -17 -113
rect 17 -147 51 -113
<< ndiode >>
rect -45 17 45 45
rect -45 -17 -17 17
rect 17 -17 45 17
rect -45 -45 45 -17
<< ndiodec >>
rect -17 -17 17 17
<< locali >>
rect -147 113 -51 147
rect -17 113 17 147
rect 51 113 147 147
rect -147 51 -113 113
rect 113 51 147 113
rect -147 -17 -113 17
rect -49 17 49 33
rect -49 -17 -17 17
rect 17 -17 49 17
rect -49 -33 49 -17
rect 113 -17 147 17
rect -147 -113 -113 -51
rect 113 -113 147 -51
rect -147 -147 -51 -113
rect -17 -147 17 -113
rect 51 -147 147 -113
<< viali >>
rect -17 -17 17 17
<< metal1 >>
rect -45 17 45 39
rect -45 -17 -17 17
rect 17 -17 45 17
rect -45 -39 45 -17
<< properties >>
string FIXED_BBOX -130 -130 130 130
<< end >>
