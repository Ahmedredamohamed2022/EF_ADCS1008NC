magic
tech sky130A
magscale 1 2
timestamp 1699926577
<< nwell >>
rect 301 1424 2543 1830
rect 301 482 616 1424
rect 2228 482 2543 1424
rect 301 373 2543 482
rect 301 -1994 616 373
rect 1957 -297 2543 373
rect 2228 -1994 2543 -297
rect 301 -2311 2543 -1994
<< mvnsubdiff >>
rect 367 1744 2477 1764
rect 367 1710 453 1744
rect 487 1710 521 1744
rect 555 1710 589 1744
rect 623 1710 657 1744
rect 691 1710 725 1744
rect 759 1710 793 1744
rect 827 1710 861 1744
rect 895 1710 929 1744
rect 963 1710 997 1744
rect 1031 1710 1065 1744
rect 1099 1710 1133 1744
rect 1167 1710 1201 1744
rect 1235 1710 1269 1744
rect 1303 1710 1337 1744
rect 1371 1710 1405 1744
rect 1439 1710 1473 1744
rect 1507 1710 1541 1744
rect 1575 1710 1609 1744
rect 1643 1710 1677 1744
rect 1711 1710 1745 1744
rect 1779 1710 1813 1744
rect 1847 1710 1881 1744
rect 1915 1710 1949 1744
rect 1983 1710 2017 1744
rect 2051 1710 2085 1744
rect 2119 1710 2153 1744
rect 2187 1710 2221 1744
rect 2255 1710 2289 1744
rect 2323 1710 2357 1744
rect 2391 1710 2477 1744
rect 367 1690 2477 1710
rect 367 1681 441 1690
rect 367 1647 387 1681
rect 421 1647 441 1681
rect 367 1613 441 1647
rect 367 1579 387 1613
rect 421 1579 441 1613
rect 367 1545 441 1579
rect 367 1511 387 1545
rect 421 1511 441 1545
rect 367 1477 441 1511
rect 367 1443 387 1477
rect 421 1443 441 1477
rect 367 1409 441 1443
rect 367 1375 387 1409
rect 421 1375 441 1409
rect 367 1341 441 1375
rect 367 1307 387 1341
rect 421 1307 441 1341
rect 367 1273 441 1307
rect 367 1239 387 1273
rect 421 1239 441 1273
rect 367 1205 441 1239
rect 367 1171 387 1205
rect 421 1171 441 1205
rect 367 1137 441 1171
rect 367 1103 387 1137
rect 421 1103 441 1137
rect 367 1069 441 1103
rect 367 1035 387 1069
rect 421 1035 441 1069
rect 367 1001 441 1035
rect 367 967 387 1001
rect 421 967 441 1001
rect 367 933 441 967
rect 367 899 387 933
rect 421 899 441 933
rect 367 865 441 899
rect 367 831 387 865
rect 421 831 441 865
rect 367 797 441 831
rect 367 763 387 797
rect 421 763 441 797
rect 367 729 441 763
rect 367 695 387 729
rect 421 695 441 729
rect 367 661 441 695
rect 367 627 387 661
rect 421 627 441 661
rect 367 593 441 627
rect 367 559 387 593
rect 421 559 441 593
rect 367 525 441 559
rect 367 491 387 525
rect 421 491 441 525
rect 367 457 441 491
rect 367 423 387 457
rect 421 423 441 457
rect 367 389 441 423
rect 367 355 387 389
rect 421 355 441 389
rect 367 321 441 355
rect 367 287 387 321
rect 421 287 441 321
rect 367 253 441 287
rect 367 219 387 253
rect 421 219 441 253
rect 367 185 441 219
rect 367 151 387 185
rect 421 151 441 185
rect 367 117 441 151
rect 367 83 387 117
rect 421 83 441 117
rect 367 49 441 83
rect 367 15 387 49
rect 421 15 441 49
rect 367 -19 441 15
rect 367 -53 387 -19
rect 421 -53 441 -19
rect 367 -87 441 -53
rect 367 -121 387 -87
rect 421 -121 441 -87
rect 367 -155 441 -121
rect 367 -189 387 -155
rect 421 -189 441 -155
rect 367 -223 441 -189
rect 367 -257 387 -223
rect 421 -257 441 -223
rect 367 -291 441 -257
rect 367 -325 387 -291
rect 421 -325 441 -291
rect 367 -359 441 -325
rect 367 -393 387 -359
rect 421 -393 441 -359
rect 367 -427 441 -393
rect 367 -461 387 -427
rect 421 -461 441 -427
rect 367 -495 441 -461
rect 367 -529 387 -495
rect 421 -529 441 -495
rect 367 -563 441 -529
rect 367 -597 387 -563
rect 421 -597 441 -563
rect 367 -631 441 -597
rect 367 -665 387 -631
rect 421 -665 441 -631
rect 367 -699 441 -665
rect 367 -733 387 -699
rect 421 -733 441 -699
rect 367 -767 441 -733
rect 367 -801 387 -767
rect 421 -801 441 -767
rect 367 -835 441 -801
rect 367 -869 387 -835
rect 421 -869 441 -835
rect 367 -903 441 -869
rect 367 -937 387 -903
rect 421 -937 441 -903
rect 367 -971 441 -937
rect 367 -1005 387 -971
rect 421 -1005 441 -971
rect 367 -1039 441 -1005
rect 367 -1073 387 -1039
rect 421 -1073 441 -1039
rect 367 -1107 441 -1073
rect 367 -1141 387 -1107
rect 421 -1141 441 -1107
rect 367 -1175 441 -1141
rect 367 -1209 387 -1175
rect 421 -1209 441 -1175
rect 367 -1243 441 -1209
rect 367 -1277 387 -1243
rect 421 -1277 441 -1243
rect 367 -1311 441 -1277
rect 367 -1345 387 -1311
rect 421 -1345 441 -1311
rect 367 -1379 441 -1345
rect 367 -1413 387 -1379
rect 421 -1413 441 -1379
rect 367 -1447 441 -1413
rect 367 -1481 387 -1447
rect 421 -1481 441 -1447
rect 367 -1515 441 -1481
rect 367 -1549 387 -1515
rect 421 -1549 441 -1515
rect 367 -1583 441 -1549
rect 367 -1617 387 -1583
rect 421 -1617 441 -1583
rect 367 -1651 441 -1617
rect 367 -1685 387 -1651
rect 421 -1685 441 -1651
rect 367 -1719 441 -1685
rect 367 -1753 387 -1719
rect 421 -1753 441 -1719
rect 367 -1787 441 -1753
rect 367 -1821 387 -1787
rect 421 -1821 441 -1787
rect 367 -1855 441 -1821
rect 367 -1889 387 -1855
rect 421 -1889 441 -1855
rect 367 -1923 441 -1889
rect 367 -1957 387 -1923
rect 421 -1957 441 -1923
rect 367 -1991 441 -1957
rect 367 -2025 387 -1991
rect 421 -2025 441 -1991
rect 367 -2059 441 -2025
rect 367 -2093 387 -2059
rect 421 -2093 441 -2059
rect 367 -2127 441 -2093
rect 367 -2161 387 -2127
rect 421 -2161 441 -2127
rect 367 -2169 441 -2161
rect 2403 1681 2477 1690
rect 2403 1647 2423 1681
rect 2457 1647 2477 1681
rect 2403 1613 2477 1647
rect 2403 1579 2423 1613
rect 2457 1579 2477 1613
rect 2403 1545 2477 1579
rect 2403 1511 2423 1545
rect 2457 1511 2477 1545
rect 2403 1477 2477 1511
rect 2403 1443 2423 1477
rect 2457 1443 2477 1477
rect 2403 1409 2477 1443
rect 2403 1375 2423 1409
rect 2457 1375 2477 1409
rect 2403 1341 2477 1375
rect 2403 1307 2423 1341
rect 2457 1307 2477 1341
rect 2403 1273 2477 1307
rect 2403 1239 2423 1273
rect 2457 1239 2477 1273
rect 2403 1205 2477 1239
rect 2403 1171 2423 1205
rect 2457 1171 2477 1205
rect 2403 1137 2477 1171
rect 2403 1103 2423 1137
rect 2457 1103 2477 1137
rect 2403 1069 2477 1103
rect 2403 1035 2423 1069
rect 2457 1035 2477 1069
rect 2403 1001 2477 1035
rect 2403 967 2423 1001
rect 2457 967 2477 1001
rect 2403 933 2477 967
rect 2403 899 2423 933
rect 2457 899 2477 933
rect 2403 865 2477 899
rect 2403 831 2423 865
rect 2457 831 2477 865
rect 2403 797 2477 831
rect 2403 763 2423 797
rect 2457 763 2477 797
rect 2403 729 2477 763
rect 2403 695 2423 729
rect 2457 695 2477 729
rect 2403 661 2477 695
rect 2403 627 2423 661
rect 2457 627 2477 661
rect 2403 593 2477 627
rect 2403 559 2423 593
rect 2457 559 2477 593
rect 2403 525 2477 559
rect 2403 491 2423 525
rect 2457 491 2477 525
rect 2403 457 2477 491
rect 2403 423 2423 457
rect 2457 423 2477 457
rect 2403 389 2477 423
rect 2403 355 2423 389
rect 2457 355 2477 389
rect 2403 321 2477 355
rect 2403 287 2423 321
rect 2457 287 2477 321
rect 2403 253 2477 287
rect 2403 219 2423 253
rect 2457 219 2477 253
rect 2403 185 2477 219
rect 2403 151 2423 185
rect 2457 151 2477 185
rect 2403 117 2477 151
rect 2403 83 2423 117
rect 2457 83 2477 117
rect 2403 49 2477 83
rect 2403 15 2423 49
rect 2457 15 2477 49
rect 2403 -19 2477 15
rect 2403 -53 2423 -19
rect 2457 -53 2477 -19
rect 2403 -87 2477 -53
rect 2403 -121 2423 -87
rect 2457 -121 2477 -87
rect 2403 -155 2477 -121
rect 2403 -189 2423 -155
rect 2457 -189 2477 -155
rect 2403 -223 2477 -189
rect 2403 -257 2423 -223
rect 2457 -257 2477 -223
rect 2403 -291 2477 -257
rect 2403 -325 2423 -291
rect 2457 -325 2477 -291
rect 2403 -359 2477 -325
rect 2403 -393 2423 -359
rect 2457 -393 2477 -359
rect 2403 -427 2477 -393
rect 2403 -461 2423 -427
rect 2457 -461 2477 -427
rect 2403 -495 2477 -461
rect 2403 -529 2423 -495
rect 2457 -529 2477 -495
rect 2403 -563 2477 -529
rect 2403 -597 2423 -563
rect 2457 -597 2477 -563
rect 2403 -631 2477 -597
rect 2403 -665 2423 -631
rect 2457 -665 2477 -631
rect 2403 -699 2477 -665
rect 2403 -733 2423 -699
rect 2457 -733 2477 -699
rect 2403 -767 2477 -733
rect 2403 -801 2423 -767
rect 2457 -801 2477 -767
rect 2403 -835 2477 -801
rect 2403 -869 2423 -835
rect 2457 -869 2477 -835
rect 2403 -903 2477 -869
rect 2403 -937 2423 -903
rect 2457 -937 2477 -903
rect 2403 -971 2477 -937
rect 2403 -1005 2423 -971
rect 2457 -1005 2477 -971
rect 2403 -1039 2477 -1005
rect 2403 -1073 2423 -1039
rect 2457 -1073 2477 -1039
rect 2403 -1107 2477 -1073
rect 2403 -1141 2423 -1107
rect 2457 -1141 2477 -1107
rect 2403 -1175 2477 -1141
rect 2403 -1209 2423 -1175
rect 2457 -1209 2477 -1175
rect 2403 -1243 2477 -1209
rect 2403 -1277 2423 -1243
rect 2457 -1277 2477 -1243
rect 2403 -1311 2477 -1277
rect 2403 -1345 2423 -1311
rect 2457 -1345 2477 -1311
rect 2403 -1379 2477 -1345
rect 2403 -1413 2423 -1379
rect 2457 -1413 2477 -1379
rect 2403 -1447 2477 -1413
rect 2403 -1481 2423 -1447
rect 2457 -1481 2477 -1447
rect 2403 -1515 2477 -1481
rect 2403 -1549 2423 -1515
rect 2457 -1549 2477 -1515
rect 2403 -1583 2477 -1549
rect 2403 -1617 2423 -1583
rect 2457 -1617 2477 -1583
rect 2403 -1651 2477 -1617
rect 2403 -1685 2423 -1651
rect 2457 -1685 2477 -1651
rect 2403 -1719 2477 -1685
rect 2403 -1753 2423 -1719
rect 2457 -1753 2477 -1719
rect 2403 -1787 2477 -1753
rect 2403 -1821 2423 -1787
rect 2457 -1821 2477 -1787
rect 2403 -1855 2477 -1821
rect 2403 -1889 2423 -1855
rect 2457 -1889 2477 -1855
rect 2403 -1923 2477 -1889
rect 2403 -1957 2423 -1923
rect 2457 -1957 2477 -1923
rect 2403 -1991 2477 -1957
rect 2403 -2025 2423 -1991
rect 2457 -2025 2477 -1991
rect 2403 -2059 2477 -2025
rect 2403 -2093 2423 -2059
rect 2457 -2093 2477 -2059
rect 2403 -2127 2477 -2093
rect 2403 -2161 2423 -2127
rect 2457 -2161 2477 -2127
rect 2403 -2169 2477 -2161
rect 367 -2189 2477 -2169
rect 367 -2223 453 -2189
rect 487 -2223 521 -2189
rect 555 -2223 589 -2189
rect 623 -2223 657 -2189
rect 691 -2223 725 -2189
rect 759 -2223 793 -2189
rect 827 -2223 861 -2189
rect 895 -2223 929 -2189
rect 963 -2223 997 -2189
rect 1031 -2223 1065 -2189
rect 1099 -2223 1133 -2189
rect 1167 -2223 1201 -2189
rect 1235 -2223 1269 -2189
rect 1303 -2223 1337 -2189
rect 1371 -2223 1405 -2189
rect 1439 -2223 1473 -2189
rect 1507 -2223 1541 -2189
rect 1575 -2223 1609 -2189
rect 1643 -2223 1677 -2189
rect 1711 -2223 1745 -2189
rect 1779 -2223 1813 -2189
rect 1847 -2223 1881 -2189
rect 1915 -2223 1949 -2189
rect 1983 -2223 2017 -2189
rect 2051 -2223 2085 -2189
rect 2119 -2223 2153 -2189
rect 2187 -2223 2221 -2189
rect 2255 -2223 2289 -2189
rect 2323 -2223 2357 -2189
rect 2391 -2223 2477 -2189
rect 367 -2243 2477 -2223
<< mvnsubdiffcont >>
rect 453 1710 487 1744
rect 521 1710 555 1744
rect 589 1710 623 1744
rect 657 1710 691 1744
rect 725 1710 759 1744
rect 793 1710 827 1744
rect 861 1710 895 1744
rect 929 1710 963 1744
rect 997 1710 1031 1744
rect 1065 1710 1099 1744
rect 1133 1710 1167 1744
rect 1201 1710 1235 1744
rect 1269 1710 1303 1744
rect 1337 1710 1371 1744
rect 1405 1710 1439 1744
rect 1473 1710 1507 1744
rect 1541 1710 1575 1744
rect 1609 1710 1643 1744
rect 1677 1710 1711 1744
rect 1745 1710 1779 1744
rect 1813 1710 1847 1744
rect 1881 1710 1915 1744
rect 1949 1710 1983 1744
rect 2017 1710 2051 1744
rect 2085 1710 2119 1744
rect 2153 1710 2187 1744
rect 2221 1710 2255 1744
rect 2289 1710 2323 1744
rect 2357 1710 2391 1744
rect 387 1647 421 1681
rect 387 1579 421 1613
rect 387 1511 421 1545
rect 387 1443 421 1477
rect 387 1375 421 1409
rect 387 1307 421 1341
rect 387 1239 421 1273
rect 387 1171 421 1205
rect 387 1103 421 1137
rect 387 1035 421 1069
rect 387 967 421 1001
rect 387 899 421 933
rect 387 831 421 865
rect 387 763 421 797
rect 387 695 421 729
rect 387 627 421 661
rect 387 559 421 593
rect 387 491 421 525
rect 387 423 421 457
rect 387 355 421 389
rect 387 287 421 321
rect 387 219 421 253
rect 387 151 421 185
rect 387 83 421 117
rect 387 15 421 49
rect 387 -53 421 -19
rect 387 -121 421 -87
rect 387 -189 421 -155
rect 387 -257 421 -223
rect 387 -325 421 -291
rect 387 -393 421 -359
rect 387 -461 421 -427
rect 387 -529 421 -495
rect 387 -597 421 -563
rect 387 -665 421 -631
rect 387 -733 421 -699
rect 387 -801 421 -767
rect 387 -869 421 -835
rect 387 -937 421 -903
rect 387 -1005 421 -971
rect 387 -1073 421 -1039
rect 387 -1141 421 -1107
rect 387 -1209 421 -1175
rect 387 -1277 421 -1243
rect 387 -1345 421 -1311
rect 387 -1413 421 -1379
rect 387 -1481 421 -1447
rect 387 -1549 421 -1515
rect 387 -1617 421 -1583
rect 387 -1685 421 -1651
rect 387 -1753 421 -1719
rect 387 -1821 421 -1787
rect 387 -1889 421 -1855
rect 387 -1957 421 -1923
rect 387 -2025 421 -1991
rect 387 -2093 421 -2059
rect 387 -2161 421 -2127
rect 2423 1647 2457 1681
rect 2423 1579 2457 1613
rect 2423 1511 2457 1545
rect 2423 1443 2457 1477
rect 2423 1375 2457 1409
rect 2423 1307 2457 1341
rect 2423 1239 2457 1273
rect 2423 1171 2457 1205
rect 2423 1103 2457 1137
rect 2423 1035 2457 1069
rect 2423 967 2457 1001
rect 2423 899 2457 933
rect 2423 831 2457 865
rect 2423 763 2457 797
rect 2423 695 2457 729
rect 2423 627 2457 661
rect 2423 559 2457 593
rect 2423 491 2457 525
rect 2423 423 2457 457
rect 2423 355 2457 389
rect 2423 287 2457 321
rect 2423 219 2457 253
rect 2423 151 2457 185
rect 2423 83 2457 117
rect 2423 15 2457 49
rect 2423 -53 2457 -19
rect 2423 -121 2457 -87
rect 2423 -189 2457 -155
rect 2423 -257 2457 -223
rect 2423 -325 2457 -291
rect 2423 -393 2457 -359
rect 2423 -461 2457 -427
rect 2423 -529 2457 -495
rect 2423 -597 2457 -563
rect 2423 -665 2457 -631
rect 2423 -733 2457 -699
rect 2423 -801 2457 -767
rect 2423 -869 2457 -835
rect 2423 -937 2457 -903
rect 2423 -1005 2457 -971
rect 2423 -1073 2457 -1039
rect 2423 -1141 2457 -1107
rect 2423 -1209 2457 -1175
rect 2423 -1277 2457 -1243
rect 2423 -1345 2457 -1311
rect 2423 -1413 2457 -1379
rect 2423 -1481 2457 -1447
rect 2423 -1549 2457 -1515
rect 2423 -1617 2457 -1583
rect 2423 -1685 2457 -1651
rect 2423 -1753 2457 -1719
rect 2423 -1821 2457 -1787
rect 2423 -1889 2457 -1855
rect 2423 -1957 2457 -1923
rect 2423 -2025 2457 -1991
rect 2423 -2093 2457 -2059
rect 2423 -2161 2457 -2127
rect 453 -2223 487 -2189
rect 521 -2223 555 -2189
rect 589 -2223 623 -2189
rect 657 -2223 691 -2189
rect 725 -2223 759 -2189
rect 793 -2223 827 -2189
rect 861 -2223 895 -2189
rect 929 -2223 963 -2189
rect 997 -2223 1031 -2189
rect 1065 -2223 1099 -2189
rect 1133 -2223 1167 -2189
rect 1201 -2223 1235 -2189
rect 1269 -2223 1303 -2189
rect 1337 -2223 1371 -2189
rect 1405 -2223 1439 -2189
rect 1473 -2223 1507 -2189
rect 1541 -2223 1575 -2189
rect 1609 -2223 1643 -2189
rect 1677 -2223 1711 -2189
rect 1745 -2223 1779 -2189
rect 1813 -2223 1847 -2189
rect 1881 -2223 1915 -2189
rect 1949 -2223 1983 -2189
rect 2017 -2223 2051 -2189
rect 2085 -2223 2119 -2189
rect 2153 -2223 2187 -2189
rect 2221 -2223 2255 -2189
rect 2289 -2223 2323 -2189
rect 2357 -2223 2391 -2189
<< locali >>
rect 387 1710 453 1744
rect 487 1710 521 1744
rect 555 1710 589 1744
rect 623 1710 657 1744
rect 691 1710 725 1744
rect 759 1710 793 1744
rect 827 1710 861 1744
rect 895 1710 929 1744
rect 963 1710 997 1744
rect 1031 1710 1065 1744
rect 1099 1710 1133 1744
rect 1167 1710 1201 1744
rect 1235 1710 1269 1744
rect 1303 1710 1337 1744
rect 1371 1710 1405 1744
rect 1439 1710 1473 1744
rect 1507 1710 1541 1744
rect 1575 1710 1609 1744
rect 1643 1710 1677 1744
rect 1711 1710 1745 1744
rect 1779 1710 1813 1744
rect 1847 1710 1881 1744
rect 1915 1710 1949 1744
rect 1983 1710 2017 1744
rect 2051 1710 2085 1744
rect 2119 1710 2153 1744
rect 2187 1710 2221 1744
rect 2255 1710 2289 1744
rect 2323 1710 2357 1744
rect 2391 1710 2457 1744
rect 387 1681 2457 1710
rect 421 1647 2423 1681
rect 387 1621 2457 1647
rect 387 1613 571 1621
rect 421 1579 571 1613
rect 387 1545 571 1579
rect 421 1511 571 1545
rect 387 1477 571 1511
rect 421 1443 571 1477
rect 387 1409 571 1443
rect 421 1375 571 1409
rect 2325 1613 2457 1621
rect 2325 1579 2423 1613
rect 2325 1545 2457 1579
rect 2325 1511 2423 1545
rect 2325 1477 2457 1511
rect 2325 1443 2423 1477
rect 2325 1409 2457 1443
rect 387 1341 571 1375
rect 421 1307 571 1341
rect 387 1273 571 1307
rect 421 1239 571 1273
rect 387 1205 571 1239
rect 421 1171 571 1205
rect 387 1137 571 1171
rect 421 1103 571 1137
rect 387 1069 571 1103
rect 421 1035 571 1069
rect 387 1001 571 1035
rect 421 967 571 1001
rect 387 933 571 967
rect 421 899 571 933
rect 387 865 571 899
rect 421 831 571 865
rect 387 797 571 831
rect 421 763 571 797
rect 387 729 571 763
rect 421 695 571 729
rect 387 661 571 695
rect 421 627 571 661
rect 387 593 571 627
rect 421 559 571 593
rect 387 525 571 559
rect 616 556 768 1376
rect 1169 1319 1343 1377
rect 1169 1285 1242 1319
rect 1276 1285 1343 1319
rect 1169 1247 1343 1285
rect 1169 1213 1242 1247
rect 1276 1213 1343 1247
rect 1169 1175 1343 1213
rect 1169 1141 1242 1175
rect 1276 1141 1343 1175
rect 1169 1103 1343 1141
rect 1169 1069 1242 1103
rect 1276 1069 1343 1103
rect 1169 1031 1343 1069
rect 1169 997 1242 1031
rect 1276 997 1343 1031
rect 1169 959 1343 997
rect 1169 925 1242 959
rect 1276 925 1343 959
rect 1169 887 1343 925
rect 1169 853 1242 887
rect 1276 853 1343 887
rect 1169 815 1343 853
rect 1169 781 1242 815
rect 1276 781 1343 815
rect 1169 743 1343 781
rect 1169 709 1242 743
rect 1276 709 1343 743
rect 1169 556 1343 709
rect 1753 1321 2255 1377
rect 1753 1287 1823 1321
rect 1857 1287 2255 1321
rect 1753 1249 2255 1287
rect 1753 1215 1823 1249
rect 1857 1215 2255 1249
rect 1753 1177 2255 1215
rect 1753 1143 1823 1177
rect 1857 1143 2255 1177
rect 1753 1105 2255 1143
rect 1753 1071 1823 1105
rect 1857 1071 2255 1105
rect 1753 1033 2255 1071
rect 1753 999 1823 1033
rect 1857 999 2255 1033
rect 1753 961 2255 999
rect 1753 927 1823 961
rect 1857 927 2255 961
rect 1753 889 2255 927
rect 1753 855 1823 889
rect 1857 855 2255 889
rect 1753 847 2255 855
rect 1753 817 1927 847
rect 1753 783 1823 817
rect 1857 783 1927 817
rect 1753 745 1927 783
rect 1753 711 1823 745
rect 1857 711 1927 745
rect 1753 556 1927 711
rect 2164 556 2255 847
rect 2325 1375 2423 1409
rect 2325 1341 2457 1375
rect 2325 1307 2423 1341
rect 2325 1273 2457 1307
rect 2325 1239 2423 1273
rect 2325 1205 2457 1239
rect 2325 1171 2423 1205
rect 2325 1137 2457 1171
rect 2325 1103 2423 1137
rect 2325 1069 2457 1103
rect 2325 1035 2423 1069
rect 2325 1001 2457 1035
rect 2325 967 2423 1001
rect 2325 933 2457 967
rect 2325 899 2423 933
rect 2325 865 2457 899
rect 2325 831 2423 865
rect 2325 797 2457 831
rect 2325 763 2423 797
rect 2325 729 2457 763
rect 2325 695 2423 729
rect 2325 661 2457 695
rect 2325 627 2423 661
rect 2325 593 2457 627
rect 2325 559 2423 593
rect 421 491 571 525
rect 387 482 571 491
rect 2325 525 2457 559
rect 2325 491 2423 525
rect 2325 482 2457 491
rect 387 457 2457 482
rect 421 423 2423 457
rect 387 389 2457 423
rect 421 355 2423 389
rect 387 342 2457 355
rect 387 321 712 342
rect 421 287 712 321
rect 387 253 712 287
rect 421 219 712 253
rect 387 185 712 219
rect 421 151 712 185
rect 387 117 712 151
rect 421 83 712 117
rect 387 49 712 83
rect 421 15 712 49
rect 387 -19 712 15
rect 421 -53 712 -19
rect 387 -87 712 -53
rect 421 -121 712 -87
rect 387 -155 712 -121
rect 421 -158 712 -155
rect 1870 321 2457 342
rect 1870 287 2423 321
rect 1870 253 2457 287
rect 1870 219 2423 253
rect 1870 185 2457 219
rect 1870 151 2423 185
rect 1870 117 2457 151
rect 1870 83 2423 117
rect 1870 49 2457 83
rect 1870 15 2423 49
rect 1870 -19 2457 15
rect 1870 -53 2423 -19
rect 1870 -87 2457 -53
rect 1870 -121 2423 -87
rect 1870 -155 2457 -121
rect 1870 -158 2423 -155
rect 421 -189 2423 -158
rect 387 -219 2457 -189
rect 387 -223 556 -219
rect 421 -257 556 -223
rect 387 -291 556 -257
rect 421 -325 556 -291
rect 2318 -223 2457 -219
rect 2318 -257 2423 -223
rect 2318 -291 2457 -257
rect 2318 -325 2423 -291
rect 387 -359 2457 -325
rect 421 -374 2423 -359
rect 421 -393 712 -374
rect 387 -427 712 -393
rect 421 -461 712 -427
rect 387 -495 712 -461
rect 421 -529 712 -495
rect 387 -563 712 -529
rect 421 -597 712 -563
rect 387 -631 712 -597
rect 421 -665 712 -631
rect 387 -699 712 -665
rect 421 -733 712 -699
rect 387 -767 712 -733
rect 421 -801 712 -767
rect 387 -835 712 -801
rect 421 -869 712 -835
rect 387 -894 712 -869
rect 2140 -393 2423 -374
rect 2140 -427 2457 -393
rect 2140 -461 2423 -427
rect 2140 -495 2457 -461
rect 2140 -529 2423 -495
rect 2140 -563 2457 -529
rect 2140 -597 2423 -563
rect 2140 -631 2457 -597
rect 2140 -665 2423 -631
rect 2140 -699 2457 -665
rect 2140 -733 2423 -699
rect 2140 -767 2457 -733
rect 2140 -801 2423 -767
rect 2140 -835 2457 -801
rect 2140 -869 2423 -835
rect 2140 -894 2457 -869
rect 387 -903 2457 -894
rect 421 -937 2423 -903
rect 387 -971 2457 -937
rect 421 -988 2423 -971
rect 421 -1005 528 -988
rect 387 -1039 528 -1005
rect 421 -1073 528 -1039
rect 2302 -1005 2423 -988
rect 2302 -1039 2457 -1005
rect 387 -1107 528 -1073
rect 421 -1141 528 -1107
rect 387 -1175 528 -1141
rect 421 -1209 528 -1175
rect 387 -1243 528 -1209
rect 421 -1277 528 -1243
rect 387 -1311 528 -1277
rect 421 -1345 528 -1311
rect 387 -1379 528 -1345
rect 421 -1413 528 -1379
rect 387 -1447 528 -1413
rect 421 -1481 528 -1447
rect 387 -1515 528 -1481
rect 421 -1549 528 -1515
rect 387 -1583 528 -1549
rect 421 -1617 528 -1583
rect 387 -1651 528 -1617
rect 421 -1685 528 -1651
rect 387 -1719 528 -1685
rect 421 -1753 528 -1719
rect 387 -1787 528 -1753
rect 421 -1821 528 -1787
rect 387 -1828 528 -1821
rect 599 -1155 2235 -1066
rect 387 -1855 421 -1828
rect 599 -1870 714 -1155
rect 2120 -1870 2235 -1155
rect 2302 -1073 2423 -1039
rect 2302 -1107 2457 -1073
rect 2302 -1141 2423 -1107
rect 2302 -1175 2457 -1141
rect 2302 -1209 2423 -1175
rect 2302 -1243 2457 -1209
rect 2302 -1277 2423 -1243
rect 2302 -1311 2457 -1277
rect 2302 -1345 2423 -1311
rect 2302 -1379 2457 -1345
rect 2302 -1413 2423 -1379
rect 2302 -1447 2457 -1413
rect 2302 -1481 2423 -1447
rect 2302 -1515 2457 -1481
rect 2302 -1549 2423 -1515
rect 2302 -1583 2457 -1549
rect 2302 -1617 2423 -1583
rect 2302 -1651 2457 -1617
rect 2302 -1685 2423 -1651
rect 2302 -1719 2457 -1685
rect 2302 -1753 2423 -1719
rect 2302 -1787 2457 -1753
rect 2302 -1821 2423 -1787
rect 2423 -1855 2457 -1821
rect 387 -1923 421 -1889
rect 387 -1991 421 -1957
rect 387 -2059 421 -2025
rect 387 -2127 421 -2093
rect 471 -1943 2378 -1870
rect 471 -2049 609 -1943
rect 2299 -2049 2378 -1943
rect 471 -2143 2378 -2049
rect 2423 -1923 2457 -1889
rect 2423 -1991 2457 -1957
rect 2423 -2059 2457 -2025
rect 2423 -2127 2457 -2093
rect 387 -2189 421 -2161
rect 2423 -2189 2457 -2161
rect 387 -2223 453 -2189
rect 487 -2223 521 -2189
rect 555 -2223 589 -2189
rect 623 -2223 657 -2189
rect 691 -2223 725 -2189
rect 759 -2223 793 -2189
rect 827 -2223 861 -2189
rect 895 -2223 929 -2189
rect 963 -2223 997 -2189
rect 1031 -2223 1065 -2189
rect 1099 -2223 1133 -2189
rect 1167 -2223 1201 -2189
rect 1235 -2223 1269 -2189
rect 1303 -2223 1337 -2189
rect 1371 -2223 1405 -2189
rect 1439 -2223 1473 -2189
rect 1507 -2223 1541 -2189
rect 1575 -2223 1609 -2189
rect 1643 -2223 1677 -2189
rect 1711 -2223 1745 -2189
rect 1779 -2223 1813 -2189
rect 1847 -2223 1881 -2189
rect 1915 -2223 1949 -2189
rect 1983 -2223 2017 -2189
rect 2051 -2223 2085 -2189
rect 2119 -2223 2153 -2189
rect 2187 -2223 2221 -2189
rect 2255 -2223 2289 -2189
rect 2323 -2223 2357 -2189
rect 2391 -2223 2457 -2189
<< viali >>
rect 1242 1285 1276 1319
rect 1242 1213 1276 1247
rect 1242 1141 1276 1175
rect 1242 1069 1276 1103
rect 1242 997 1276 1031
rect 1242 925 1276 959
rect 1242 853 1276 887
rect 1242 781 1276 815
rect 1242 709 1276 743
rect 1823 1287 1857 1321
rect 1823 1215 1857 1249
rect 1823 1143 1857 1177
rect 1823 1071 1857 1105
rect 1823 999 1857 1033
rect 1823 927 1857 961
rect 1823 855 1857 889
rect 1823 783 1857 817
rect 1823 711 1857 745
rect 556 -325 2318 -219
rect 609 -2049 2299 -1943
<< metal1 >>
rect 393 1521 2463 1563
rect 393 1341 571 1521
rect 815 1341 2463 1521
rect 393 1321 2463 1341
rect 393 1319 1823 1321
rect 393 1306 1242 1319
rect 824 764 888 1306
rect 1211 1285 1242 1306
rect 1276 1306 1823 1319
rect 1276 1285 1308 1306
rect 1211 1247 1308 1285
rect 340 619 540 690
rect 943 619 980 1231
rect 1211 1213 1242 1247
rect 1276 1213 1308 1247
rect 1211 1175 1308 1213
rect 340 567 907 619
rect 959 567 980 619
rect 340 490 540 567
rect 943 401 980 567
rect 1052 502 1101 1172
rect 1211 1141 1242 1175
rect 1276 1141 1308 1175
rect 1211 1103 1308 1141
rect 1211 1069 1242 1103
rect 1276 1069 1308 1103
rect 1211 1031 1308 1069
rect 1211 997 1242 1031
rect 1276 997 1308 1031
rect 1211 959 1308 997
rect 1211 925 1242 959
rect 1276 925 1308 959
rect 1211 887 1308 925
rect 1211 853 1242 887
rect 1276 853 1308 887
rect 1211 815 1308 853
rect 1211 781 1242 815
rect 1276 781 1308 815
rect 1211 743 1308 781
rect 1406 760 1470 1306
rect 1791 1287 1823 1306
rect 1857 1306 2463 1321
rect 1857 1287 1888 1306
rect 1791 1249 1888 1287
rect 1211 709 1242 743
rect 1276 709 1308 743
rect 1211 659 1308 709
rect 1534 502 1571 1232
rect 1791 1215 1823 1249
rect 1857 1215 1888 1249
rect 1791 1177 1888 1215
rect 1052 453 1571 502
rect 909 364 1099 401
rect 909 200 946 364
rect 1062 200 1099 364
rect 793 136 866 153
rect 793 84 804 136
rect 856 84 866 136
rect 793 72 866 84
rect 793 20 804 72
rect 856 20 866 72
rect 793 8 866 20
rect 793 -44 804 8
rect 856 -44 866 8
rect 793 -59 866 -44
rect 964 -92 1036 156
rect 1158 139 1207 453
rect 1534 401 1571 453
rect 1620 500 1669 1171
rect 1791 1143 1823 1177
rect 1857 1143 1888 1177
rect 1791 1105 1888 1143
rect 1791 1071 1823 1105
rect 1857 1071 1888 1105
rect 1791 1033 1888 1071
rect 1791 999 1823 1033
rect 1857 999 1888 1033
rect 1791 961 1888 999
rect 1791 927 1823 961
rect 1857 927 1888 961
rect 1791 889 1888 927
rect 1791 855 1823 889
rect 1857 855 1888 889
rect 1791 817 1888 855
rect 1791 783 1823 817
rect 1857 783 1888 817
rect 1791 745 1888 783
rect 1791 711 1823 745
rect 1857 711 1888 745
rect 1791 664 1888 711
rect 2009 619 2080 739
rect 2009 567 2018 619
rect 2070 567 2080 619
rect 2009 561 2080 567
rect 1620 451 1792 500
rect 1490 364 1680 401
rect 1490 200 1527 364
rect 1643 200 1680 364
rect 1147 137 1207 139
rect 1147 85 1148 137
rect 1200 85 1207 137
rect 1147 73 1207 85
rect 1147 21 1148 73
rect 1200 21 1207 73
rect 1147 9 1207 21
rect 1147 -43 1148 9
rect 1200 -43 1207 9
rect 1147 -45 1207 -43
rect 1158 -57 1207 -45
rect 1375 138 1448 151
rect 1375 86 1383 138
rect 1435 86 1448 138
rect 1375 74 1448 86
rect 1375 22 1383 74
rect 1435 22 1448 74
rect 1375 10 1448 22
rect 1375 -42 1383 10
rect 1435 -42 1448 10
rect 1375 -61 1448 -42
rect 1552 -92 1624 151
rect 1743 140 1792 451
rect 1732 138 1792 140
rect 1732 86 1733 138
rect 1785 86 1792 138
rect 1732 74 1792 86
rect 1732 22 1733 74
rect 1785 22 1792 74
rect 1732 10 1792 22
rect 1732 -42 1733 10
rect 1785 -42 1792 10
rect 1732 -44 1792 -42
rect 1743 -59 1792 -44
rect 326 -219 2478 -92
rect 326 -325 556 -219
rect 2318 -325 2478 -219
rect 326 -368 2478 -325
rect 904 -449 973 -397
rect 1025 -449 1046 -397
rect 904 -453 1046 -449
rect 1370 -403 1525 -402
rect 745 -643 867 -636
rect 745 -695 779 -643
rect 831 -695 867 -643
rect 745 -701 867 -695
rect 904 -867 939 -453
rect 1370 -455 1390 -403
rect 1442 -455 1525 -403
rect 1370 -458 1525 -455
rect 1190 -517 1292 -495
rect 1190 -569 1215 -517
rect 1267 -569 1292 -517
rect 1190 -591 1292 -569
rect 977 -642 1099 -635
rect 977 -694 1012 -642
rect 1064 -694 1099 -642
rect 977 -700 1099 -694
rect 1350 -655 1452 -648
rect 1350 -707 1375 -655
rect 1427 -707 1452 -655
rect 1350 -714 1452 -707
rect 1489 -749 1525 -458
rect 1562 -517 1664 -495
rect 1562 -569 1587 -517
rect 1639 -569 1664 -517
rect 1562 -591 1664 -569
rect 1755 -512 1876 -505
rect 1755 -564 1789 -512
rect 1841 -564 1876 -512
rect 1755 -570 1876 -564
rect 1988 -512 2109 -505
rect 1988 -564 2022 -512
rect 2074 -564 2109 -512
rect 1988 -570 2109 -564
rect 1334 -783 1685 -749
rect 1334 -785 1625 -783
rect 1617 -835 1625 -785
rect 1677 -835 1685 -783
rect 1617 -839 1685 -835
rect 1913 -867 1948 -760
rect 904 -915 1948 -867
rect 2209 -776 2526 -576
rect 2209 -786 2393 -776
rect 314 -974 891 -964
rect 314 -1154 752 -974
rect 868 -1154 891 -974
rect 314 -1164 891 -1154
rect 1051 -1047 1128 -1037
rect 1051 -1099 1063 -1047
rect 1115 -1099 1128 -1047
rect 1051 -1107 1128 -1099
rect 1051 -1261 1087 -1107
rect 894 -1289 1087 -1261
rect 1479 -1264 1515 -915
rect 1728 -1047 1805 -1039
rect 1728 -1099 1740 -1047
rect 1792 -1099 1805 -1047
rect 1728 -1109 1805 -1099
rect 887 -1297 1087 -1289
rect 740 -1359 856 -1342
rect 740 -1411 772 -1359
rect 824 -1411 856 -1359
rect 740 -1423 856 -1411
rect 740 -1475 772 -1423
rect 824 -1475 856 -1423
rect 740 -1491 856 -1475
rect 887 -1784 923 -1297
rect 1322 -1300 1515 -1264
rect 1756 -1262 1792 -1109
rect 2209 -1222 2244 -786
rect 2360 -1222 2393 -786
rect 2209 -1236 2393 -1222
rect 1756 -1298 1949 -1262
rect 967 -1359 1083 -1342
rect 967 -1411 999 -1359
rect 1051 -1411 1083 -1359
rect 967 -1423 1083 -1411
rect 967 -1475 999 -1423
rect 1051 -1475 1083 -1423
rect 967 -1491 1083 -1475
rect 1323 -1362 1440 -1352
rect 1323 -1414 1355 -1362
rect 1407 -1414 1440 -1362
rect 1323 -1426 1440 -1414
rect 1323 -1478 1355 -1426
rect 1407 -1478 1440 -1426
rect 1323 -1488 1440 -1478
rect 1166 -1598 1282 -1581
rect 1166 -1650 1198 -1598
rect 1250 -1650 1282 -1598
rect 1166 -1662 1282 -1650
rect 1166 -1714 1198 -1662
rect 1250 -1714 1282 -1662
rect 1166 -1730 1282 -1714
rect 1479 -1773 1515 -1300
rect 1552 -1598 1668 -1581
rect 1552 -1650 1584 -1598
rect 1636 -1650 1668 -1598
rect 1552 -1662 1668 -1650
rect 1552 -1714 1584 -1662
rect 1636 -1714 1668 -1662
rect 1552 -1730 1668 -1714
rect 1750 -1598 1866 -1581
rect 1750 -1650 1782 -1598
rect 1834 -1650 1866 -1598
rect 1750 -1662 1866 -1650
rect 1750 -1714 1782 -1662
rect 1834 -1714 1866 -1662
rect 1750 -1730 1866 -1714
rect 1347 -1809 1515 -1773
rect 1910 -1786 1946 -1298
rect 1978 -1598 2094 -1581
rect 1978 -1650 2010 -1598
rect 2062 -1650 2094 -1598
rect 1978 -1662 2094 -1650
rect 1978 -1714 2010 -1662
rect 2062 -1714 2094 -1662
rect 1978 -1730 2094 -1714
rect 328 -1899 2515 -1870
rect 328 -2079 569 -1899
rect 813 -1943 2515 -1899
rect 2299 -2049 2515 -1943
rect 813 -2079 2515 -2049
rect 328 -2105 2515 -2079
<< via1 >>
rect 571 1341 815 1521
rect 907 567 959 619
rect 804 84 856 136
rect 804 20 856 72
rect 804 -44 856 8
rect 2018 567 2070 619
rect 1148 85 1200 137
rect 1148 21 1200 73
rect 1148 -43 1200 9
rect 1383 86 1435 138
rect 1383 22 1435 74
rect 1383 -42 1435 10
rect 1733 86 1785 138
rect 1733 22 1785 74
rect 1733 -42 1785 10
rect 973 -449 1025 -397
rect 779 -695 831 -643
rect 1390 -455 1442 -403
rect 1215 -569 1267 -517
rect 1012 -694 1064 -642
rect 1375 -707 1427 -655
rect 1587 -569 1639 -517
rect 1789 -564 1841 -512
rect 2022 -564 2074 -512
rect 1625 -835 1677 -783
rect 752 -1154 868 -974
rect 1063 -1099 1115 -1047
rect 1740 -1099 1792 -1047
rect 772 -1411 824 -1359
rect 772 -1475 824 -1423
rect 2244 -1222 2360 -786
rect 999 -1411 1051 -1359
rect 999 -1475 1051 -1423
rect 1355 -1414 1407 -1362
rect 1355 -1478 1407 -1426
rect 1198 -1650 1250 -1598
rect 1198 -1714 1250 -1662
rect 1584 -1650 1636 -1598
rect 1584 -1714 1636 -1662
rect 1782 -1650 1834 -1598
rect 1782 -1714 1834 -1662
rect 2010 -1650 2062 -1598
rect 2010 -1714 2062 -1662
rect 569 -1943 813 -1899
rect 569 -2049 609 -1943
rect 609 -2049 813 -1943
rect 569 -2079 813 -2049
<< metal2 >>
rect 529 1521 867 1556
rect 529 1341 571 1521
rect 815 1341 867 1521
rect 529 1306 867 1341
rect 529 -1870 660 1306
rect 886 567 907 619
rect 959 567 2018 619
rect 2070 567 2087 619
rect 795 137 1207 141
rect 795 136 1148 137
rect 795 84 804 136
rect 856 85 1148 136
rect 1200 85 1207 137
rect 856 84 1207 85
rect 795 73 1207 84
rect 795 72 1148 73
rect 795 20 804 72
rect 856 21 1148 72
rect 1200 21 1207 73
rect 856 20 1207 21
rect 795 9 1207 20
rect 795 8 1148 9
rect 795 -44 804 8
rect 856 -43 1148 8
rect 1200 -43 1207 9
rect 856 -44 1207 -43
rect 795 -47 1207 -44
rect 1376 138 1792 142
rect 1376 86 1383 138
rect 1435 86 1733 138
rect 1785 86 1792 138
rect 1376 74 1792 86
rect 1376 22 1383 74
rect 1435 22 1733 74
rect 1785 22 1792 74
rect 1376 10 1792 22
rect 1376 -42 1383 10
rect 1435 -42 1733 10
rect 1785 -42 1792 10
rect 1376 -46 1792 -42
rect 959 -397 1040 -47
rect 959 -449 973 -397
rect 1025 -449 1040 -397
rect 959 -455 1040 -449
rect 1376 -403 1457 -46
rect 1376 -455 1390 -403
rect 1442 -455 1457 -403
rect 1376 -461 1457 -455
rect 736 -512 2393 -489
rect 736 -517 1789 -512
rect 736 -569 1215 -517
rect 1267 -569 1587 -517
rect 1639 -564 1789 -517
rect 1841 -564 2022 -512
rect 2074 -564 2393 -512
rect 1639 -569 2393 -564
rect 736 -593 2393 -569
rect 732 -642 2127 -634
rect 732 -643 1012 -642
rect 732 -695 779 -643
rect 831 -694 1012 -643
rect 1064 -655 2127 -642
rect 1064 -694 1375 -655
rect 831 -695 1375 -694
rect 732 -707 1375 -695
rect 1427 -707 2127 -655
rect 732 -738 2127 -707
rect 732 -974 891 -738
rect 732 -1154 752 -974
rect 868 -1154 891 -974
rect 1623 -783 1679 -772
rect 1623 -835 1625 -783
rect 1677 -835 1679 -783
rect 1623 -1045 1679 -835
rect 2209 -786 2393 -593
rect 1043 -1047 1816 -1045
rect 1043 -1099 1063 -1047
rect 1115 -1099 1740 -1047
rect 1792 -1099 1816 -1047
rect 1043 -1101 1816 -1099
rect 732 -1313 891 -1154
rect 2209 -1222 2244 -786
rect 2360 -1222 2393 -786
rect 732 -1359 2122 -1313
rect 732 -1411 772 -1359
rect 824 -1411 999 -1359
rect 1051 -1362 2122 -1359
rect 1051 -1411 1355 -1362
rect 732 -1414 1355 -1411
rect 1407 -1414 2122 -1362
rect 732 -1423 2122 -1414
rect 732 -1475 772 -1423
rect 824 -1475 999 -1423
rect 1051 -1426 2122 -1423
rect 1051 -1475 1355 -1426
rect 732 -1478 1355 -1475
rect 1407 -1478 2122 -1426
rect 732 -1497 2122 -1478
rect 2209 -1558 2393 -1222
rect 733 -1598 2393 -1558
rect 733 -1650 1198 -1598
rect 1250 -1650 1584 -1598
rect 1636 -1650 1782 -1598
rect 1834 -1650 2010 -1598
rect 2062 -1650 2393 -1598
rect 733 -1662 2393 -1650
rect 733 -1714 1198 -1662
rect 1250 -1714 1584 -1662
rect 1636 -1714 1782 -1662
rect 1834 -1714 2010 -1662
rect 2062 -1714 2393 -1662
rect 733 -1742 2393 -1714
rect 529 -1899 849 -1870
rect 529 -2079 569 -1899
rect 813 -2079 849 -1899
rect 529 -2105 849 -2079
use sky130_fd_pr__pfet_g5v0d10v5_U6NWY6  sky130_fd_pr__pfet_g5v0d10v5_U6NWY6_0
timestamp 1699926577
transform 1 0 922 0 1 -638
box -308 -362 308 362
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  sky130_fd_pr__pfet_g5v0d10v5_U62SY6_0
timestamp 1699926577
transform 1 0 1585 0 -1 82
box -387 -362 387 362
use sky130_fd_pr__diode_pw2nd_05v5_FT76RJ  XD1
timestamp 1699926577
transform 1 0 2045 0 -1 703
box -173 -173 173 173
use sky130_fd_pr__nfet_g5v0d10v5_EJGQFX  XM1
timestamp 1699926577
transform -1 0 1417 0 1 -1536
box -347 -448 347 448
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM3
timestamp 1699926577
transform -1 0 907 0 1 -1536
box -268 -448 268 448
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  XM4
timestamp 1699926577
transform 1 0 1427 0 1 -638
box -387 -362 387 362
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM5
timestamp 1699926577
transform 1 0 1927 0 1 -1536
box -268 -448 268 448
use sky130_fd_pr__pfet_g5v0d10v5_U6NWY6  XM6
timestamp 1699926577
transform 1 0 1932 0 1 -638
box -308 -362 308 362
use sky130_fd_pr__pfet_g5v0d10v5_U62SY6  XM7
timestamp 1699926577
transform 1 0 1001 0 -1 82
box -387 -362 387 362
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM8
timestamp 1699926577
transform 1 0 964 0 -1 966
box -268 -448 268 448
use sky130_fd_pr__nfet_g5v0d10v5_WSEQJ8  XM10
timestamp 1699926577
transform 1 0 1546 0 -1 966
box -268 -448 268 448
<< labels >>
flabel metal1 s 1271 478 1271 478 0 FreeSans 61 0 0 0 holdb
flabel metal1 s 1705 473 1705 473 0 FreeSans 61 0 0 0 holdp
flabel metal1 s 340 490 540 690 0 FreeSans 49 0 0 0 hold
port 1 nsew
flabel metal1 s 336 -2091 536 -1891 0 FreeSans 49 0 0 0 vss
port 2 nsew
flabel metal1 s 2326 -776 2526 -576 0 FreeSans 49 0 0 0 out
port 3 nsew
flabel metal1 s 314 -1164 514 -964 0 FreeSans 49 0 0 0 in
port 4 nsew
flabel metal1 s 326 -352 526 -152 0 FreeSans 49 0 0 0 vdd
port 5 nsew
<< end >>
