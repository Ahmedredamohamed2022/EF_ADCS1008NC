VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO EF_ADCS1008NC
  CLASS BLOCK ;
  FOREIGN EF_ADCS1008NC ;
  ORIGIN 15.810 4.960 ;
  SIZE 179.285 BY 490.035 ;
  PIN VSS
    ANTENNAGATEAREA 130.000000 ;
    ANTENNADIFFAREA 530.402893 ;
    PORT
      LAYER met3 ;
        RECT 96.070 346.940 97.480 348.330 ;
    END
  END VSS
  PIN VIN[0]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 124.600 483.940 125.130 484.790 ;
    END
  END VIN[0]
  PIN VIN[1]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 107.620 484.000 108.150 484.850 ;
    END
  END VIN[1]
  PIN VIN[2]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 91.120 483.860 91.650 484.710 ;
    END
  END VIN[2]
  PIN VIN[3]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 73.820 483.800 74.350 484.650 ;
    END
  END VIN[3]
  PIN VIN[4]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 57.020 483.740 57.550 484.590 ;
    END
  END VIN[4]
  PIN VIN[5]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 39.790 483.860 40.320 484.710 ;
    END
  END VIN[5]
  PIN VIN[6]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 23.160 483.860 23.690 484.710 ;
    END
  END VIN[6]
  PIN VIN[7]
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 5.950 483.920 6.480 484.770 ;
    END
  END VIN[7]
  PIN B[0]
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 162.810 449.390 163.100 449.920 ;
    END
  END B[0]
  PIN B[1]
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 162.840 447.920 163.130 448.450 ;
    END
  END B[1]
  PIN B[2]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 162.750 446.550 163.040 447.080 ;
    END
  END B[2]
  PIN CMP
    ANTENNADIFFAREA 0.492900 ;
    PORT
      LAYER met3 ;
        RECT 162.800 422.200 163.330 422.990 ;
    END
  END CMP
  PIN RST
    ANTENNAGATEAREA 0.504000 ;
    PORT
      LAYER met3 ;
        RECT 162.740 316.550 163.210 317.150 ;
    END
  END RST
  PIN DVDD
    ANTENNAGATEAREA 47.261497 ;
    ANTENNADIFFAREA 92.613647 ;
    PORT
      LAYER met3 ;
        RECT -14.580 0.790 -13.970 1.490 ;
    END
  END DVDD
  PIN DVSS
    ANTENNAGATEAREA 74.759102 ;
    ANTENNADIFFAREA 816.096802 ;
    PORT
      LAYER met3 ;
        RECT -14.890 -1.770 -14.280 -1.070 ;
    END
  END DVSS
  PIN VDD
    ANTENNAGATEAREA 100.000000 ;
    ANTENNADIFFAREA 2017.665894 ;
    PORT
      LAYER met3 ;
        RECT -14.650 -4.290 -14.040 -3.590 ;
    END
  END VDD
  PIN DATA[0]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -14.640 13.290 -14.250 13.610 ;
    END
  END DATA[0]
  PIN DATA[1]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -14.840 49.370 -14.640 49.780 ;
    END
  END DATA[1]
  PIN VL
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met3 ;
        RECT -15.160 18.320 -14.790 18.810 ;
    END
  END VL
  PIN VH
    ANTENNADIFFAREA 26.099998 ;
    PORT
      LAYER met3 ;
        RECT -15.180 16.450 -14.810 16.940 ;
    END
  END VH
  PIN DATA[2]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -14.790 83.400 -14.490 83.780 ;
    END
  END DATA[2]
  PIN DATA[3]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -14.860 118.350 -14.470 118.930 ;
    END
  END DATA[3]
  PIN DATA[4]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -14.900 152.260 -14.340 152.650 ;
    END
  END DATA[4]
  PIN DATA[5]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -14.660 184.500 -14.300 185.060 ;
    END
  END DATA[5]
  PIN DATA[6]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -14.840 219.370 -14.580 219.770 ;
    END
  END DATA[6]
  PIN DATA[7]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -15.140 251.350 -14.940 251.600 ;
    END
  END DATA[7]
  PIN DATA[8]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -14.920 281.370 -14.620 281.710 ;
    END
  END DATA[8]
  PIN DATA[9]
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met3 ;
        RECT -14.920 317.410 -14.660 317.700 ;
    END
  END DATA[9]
  PIN EN
    ANTENNAGATEAREA 1.500000 ;
    ANTENNADIFFAREA 1.080000 ;
    PORT
      LAYER met3 ;
        RECT -15.530 384.050 -15.020 384.650 ;
    END
  END EN
  PIN HOLD
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.360000 ;
    PORT
      LAYER met3 ;
        RECT -15.710 405.380 -15.380 405.660 ;
    END
  END HOLD
  OBS
      LAYER li1 ;
        RECT -8.600 7.615 161.965 469.590 ;
      LAYER met1 ;
        RECT -15.720 5.090 162.120 469.590 ;
      LAYER met2 ;
        RECT -15.720 485.050 107.340 485.075 ;
        RECT -15.720 483.640 5.670 485.050 ;
        RECT 6.760 484.990 107.340 485.050 ;
        RECT 6.760 483.640 22.880 484.990 ;
        RECT -15.720 483.580 22.880 483.640 ;
        RECT 23.970 483.580 39.510 484.990 ;
        RECT 40.600 484.930 90.840 484.990 ;
        RECT 40.600 484.870 73.540 484.930 ;
        RECT 40.600 483.580 56.740 484.870 ;
        RECT -15.720 483.460 56.740 483.580 ;
        RECT 57.830 483.520 73.540 484.870 ;
        RECT 74.630 483.580 90.840 484.930 ;
        RECT 91.930 483.720 107.340 484.990 ;
        RECT 108.430 485.070 162.765 485.075 ;
        RECT 108.430 483.720 124.320 485.070 ;
        RECT 91.930 483.660 124.320 483.720 ;
        RECT 125.410 483.660 162.765 485.070 ;
        RECT 91.930 483.580 162.765 483.660 ;
        RECT 74.630 483.520 162.765 483.580 ;
        RECT 57.830 483.460 162.765 483.520 ;
        RECT -15.720 3.010 162.765 483.460 ;
      LAYER met3 ;
        RECT -15.810 450.320 163.475 482.050 ;
        RECT -15.810 448.990 162.410 450.320 ;
        RECT -15.810 448.850 163.475 448.990 ;
        RECT -15.810 447.520 162.440 448.850 ;
        RECT -15.810 447.480 163.475 447.520 ;
        RECT -15.810 446.150 162.350 447.480 ;
        RECT 163.440 446.150 163.475 447.480 ;
        RECT -15.810 423.390 163.475 446.150 ;
        RECT -15.810 421.800 162.400 423.390 ;
        RECT -15.810 406.060 163.475 421.800 ;
        RECT -14.980 405.840 163.475 406.060 ;
        RECT -15.810 405.660 163.475 405.840 ;
        RECT -15.810 405.380 -15.710 405.660 ;
        RECT -14.980 405.380 163.475 405.660 ;
        RECT -15.810 405.250 163.475 405.380 ;
        RECT -14.980 404.980 163.475 405.250 ;
        RECT -15.810 385.050 163.475 404.980 ;
        RECT -14.620 383.650 163.475 385.050 ;
        RECT -15.810 348.730 163.475 383.650 ;
        RECT -15.810 346.540 95.670 348.730 ;
        RECT 97.880 346.540 163.475 348.730 ;
        RECT -15.810 318.100 163.475 346.540 ;
        RECT -15.810 317.010 -15.320 318.100 ;
        RECT -14.260 317.550 163.475 318.100 ;
        RECT -14.260 317.010 162.340 317.550 ;
        RECT -15.810 316.150 162.340 317.010 ;
        RECT -15.810 282.110 163.475 316.150 ;
        RECT -15.810 280.970 -15.320 282.110 ;
        RECT -14.220 280.970 163.475 282.110 ;
        RECT -15.810 252.000 163.475 280.970 ;
        RECT -15.810 250.950 -15.540 252.000 ;
        RECT -14.540 250.950 163.475 252.000 ;
        RECT -15.810 220.170 163.475 250.950 ;
        RECT -15.810 218.970 -15.240 220.170 ;
        RECT -14.180 218.970 163.475 220.170 ;
        RECT -15.810 185.460 163.475 218.970 ;
        RECT -15.810 184.100 -15.060 185.460 ;
        RECT -13.900 184.100 163.475 185.460 ;
        RECT -15.810 153.050 163.475 184.100 ;
        RECT -15.810 151.860 -15.300 153.050 ;
        RECT -13.940 151.860 163.475 153.050 ;
        RECT -15.810 119.330 163.475 151.860 ;
        RECT -15.810 117.950 -15.260 119.330 ;
        RECT -14.070 117.950 163.475 119.330 ;
        RECT -15.810 84.180 163.475 117.950 ;
        RECT -15.810 83.000 -15.190 84.180 ;
        RECT -14.090 83.000 163.475 84.180 ;
        RECT -15.810 50.180 163.475 83.000 ;
        RECT -15.810 48.970 -15.240 50.180 ;
        RECT -14.240 48.970 163.475 50.180 ;
        RECT -15.810 19.210 163.475 48.970 ;
        RECT -15.810 17.920 -15.560 19.210 ;
        RECT -14.390 17.920 163.475 19.210 ;
        RECT -15.810 17.340 163.475 17.920 ;
        RECT -15.810 16.050 -15.580 17.340 ;
        RECT -14.410 16.050 163.475 17.340 ;
        RECT -15.810 14.010 163.475 16.050 ;
        RECT -15.810 12.890 -15.040 14.010 ;
        RECT -13.850 12.890 163.475 14.010 ;
        RECT -15.810 1.890 163.475 12.890 ;
        RECT -15.810 0.390 -14.980 1.890 ;
        RECT -13.570 0.390 163.475 1.890 ;
        RECT -15.810 -0.670 163.475 0.390 ;
        RECT -15.810 -2.170 -15.290 -0.670 ;
        RECT -13.880 -2.170 163.475 -0.670 ;
        RECT -15.810 -3.190 163.475 -2.170 ;
        RECT -15.810 -4.690 -15.050 -3.190 ;
        RECT -13.640 -4.690 163.475 -3.190 ;
        RECT -15.810 -4.860 163.475 -4.690 ;
      LAYER met4 ;
        RECT -15.140 -4.960 163.345 482.040 ;
      LAYER met5 ;
        RECT 7.815 141.020 158.600 469.590 ;
  END
END EF_ADCS1008NC
END LIBRARY

